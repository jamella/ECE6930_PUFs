
//^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^
// GF(6)
//^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^

function[11:0] fn_bch_dec_gf6;
input[62:0] d;

reg [11:0] p;
begin

 p[0] = d[0]^ d[2]^ d[6]^ d[7]^ d[9]^ d[11]^ d[12]^ d[13]^ d[16]^ d[19]^ d[22]^ d[23]^
              d[24]^ d[25]^ d[26]^ d[27]^ d[29]^ d[30]^ d[34]^ d[35]^ d[39]^ d[41]^ d[42]^ d[45]^
              d[46]^ d[47]^ d[48]^ d[51];

 p[1] = d[1]^ d[3]^ d[7]^ d[8]^ d[10]^ d[12]^ d[13]^ d[14]^ d[17]^ d[20]^ d[23]^ d[24]^
              d[25]^ d[26]^ d[27]^ d[28]^ d[30]^ d[31]^ d[35]^ d[36]^ d[40]^ d[42]^ d[43]^
              d[46]^ d[47]^ d[48]^ d[49]^ d[52];

 p[2] = d[2]^ d[4]^ d[8]^ d[9]^ d[11]^ d[13]^ d[14]^ d[15]^ d[18]^ d[21]^ d[24]^ d[25]^
              d[26]^ d[27]^ d[28]^ d[29]^ d[31]^ d[32]^ d[36]^ d[37]^ d[41]^ d[43]^ d[44]^
              d[47]^ d[48]^ d[49]^ d[50]^ d[53];

 p[3] = d[0]^ d[2]^ d[3]^ d[5]^ d[6]^ d[7]^ d[10]^ d[11]^ d[13]^ d[14]^ d[15]^ d[23]^
              d[24]^ d[28]^ d[32]^ d[33]^ d[34]^ d[35]^ d[37]^ d[38]^ d[39]^ d[41]^ d[44]^
              d[46]^ d[47]^ d[49]^ d[50]^ d[54];

 p[4] = d[0]^ d[1]^ d[2]^ d[3]^ d[4]^ d[8]^ d[9]^ d[13]^ d[14]^ d[15]^ d[19]^ d[22]^ d[23]^
              d[26]^ d[27]^ d[30]^ d[33]^ d[36]^ d[38]^ d[40]^ d[41]^ d[46]^ d[50]^ d[55];

 p[5] = d[0]^ d[1]^ d[3]^ d[4]^ d[5]^ d[6]^ d[7]^ d[10]^ d[11]^ d[12]^ d[13]^ d[14]^ d[15]^
              d[19]^ d[20]^ d[22]^ d[25]^ d[26]^ d[28]^ d[29]^ d[30]^ d[31]^ d[35]^ d[37]^ d[45]^
              d[46]^ d[48]^ d[56];

 p[6] = d[1]^ d[2]^ d[4]^ d[5]^ d[6]^ d[7]^ d[8]^ d[11]^ d[12]^ d[13]^ d[14]^ d[15]^ d[16]^
              d[20]^ d[21]^ d[23]^ d[26]^ d[27]^ d[29]^ d[30]^ d[31]^ d[32]^ d[36]^ d[38]^ d[46]^
              d[47]^ d[49]^ d[57];

 p[7] = d[2]^ d[3]^ d[5]^ d[6]^ d[7]^ d[8]^ d[9]^ d[12]^ d[13]^ d[14]^ d[15]^ d[16]^ d[17]^
              d[21]^ d[22]^ d[24]^ d[27]^ d[28]^ d[30]^ d[31]^ d[32]^ d[33]^ d[37]^ d[39]^ d[47]^
              d[48]^ d[50]^ d[58];

 p[8] = d[0]^ d[2]^ d[3]^ d[4]^ d[8]^ d[10]^ d[11]^ d[12]^ d[14]^ d[15]^ d[17]^ d[18]^ d[19]^
              d[24]^ d[26]^ d[27]^ d[28]^ d[30]^ d[31]^ d[32]^ d[33]^ d[35]^ d[38]^ d[39]^ d[40]^
              d[41]^ d[42]^ d[45]^ d[46]^ d[47]^ d[49]^ d[59];

 p[9] = d[1]^ d[3]^ d[4]^ d[5]^ d[9]^ d[11]^ d[12]^ d[13]^ d[15]^ d[16]^ d[18]^ d[19]^ d[20]^
              d[25]^ d[27]^ d[28]^ d[29]^ d[31]^ d[32]^ d[33]^ d[34]^ d[36]^ d[39]^ d[40]^ d[41]^
              d[42]^ d[43]^ d[46]^ d[47]^ d[48]^ d[50]^ d[60];

 p[10] = d[0]^ d[4]^ d[5]^ d[7]^ d[9]^ d[10]^ d[11]^ d[14]^ d[17]^ d[20]^ d[21]^ d[22]^ d[23]^
               d[24]^ d[25]^ d[27]^ d[28]^ d[32]^ d[33]^ d[37]^ d[39]^ d[40]^ d[43]^ d[44]^ d[45]^ d[46]^
               d[49]^ d[61];

 p[11] = d[1]^ d[5]^ d[6]^ d[8]^ d[10]^ d[11]^ d[12]^ d[15]^ d[18]^ d[21]^ d[22]^ d[23]^ d[24]^
               d[25]^ d[26]^ d[28]^ d[29]^ d[33]^ d[34]^ d[38]^ d[40]^ d[41]^ d[44]^ d[45]^ d[46]^ d[47]^
               d[50]^ d[62];

fn_bch_dec_gf6 = p;
end	

endfunction // fn_bch_dec_gf6

