
//&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&
// GF(6) Error pattern ROM
//&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&

function[62:0] fn_err_pat_dcd_gf6_rom;						
input[11:0]           syndromes; 

reg[62:0]            errs;   
begin
 case(syndromes)  

    12'h539 : errs =          63'b000000000000000000000000000000000000000000000000000000000000001; // S (0x0000000000000001) 
//    12'hf4b : errs =          63'b000000000000000000000000000000000000000000000000000000000000011; // D (0x0000000000000003) 
//    12'h4e4 : errs =          63'b000000000000000000000000000000000000000000000000000000000000101; // D (0x0000000000000005) 
//    12'h683 : errs =          63'b000000000000000000000000000000000000000000000000000000000001001; // D (0x0000000000000009) 
//    12'h24d : errs =          63'b000000000000000000000000000000000000000000000000000000000010001; // D (0x0000000000000011) 
//    12'hbd1 : errs =          63'b000000000000000000000000000000000000000000000000000000000100001; // D (0x0000000000000021) 
//    12'hdd0 : errs =          63'b000000000000000000000000000000000000000000000000000000001000001; // D (0x0000000000000041) 
//    12'h1d2 : errs =          63'b000000000000000000000000000000000000000000000000000000010000001; // D (0x0000000000000081) 
//    12'hcef : errs =          63'b000000000000000000000000000000000000000000000000000000100000001; // D (0x0000000000000101) 
//    12'h3ac : errs =          63'b000000000000000000000000000000000000000000000000000001000000001; // D (0x0000000000000201) 
//    12'h813 : errs =          63'b000000000000000000000000000000000000000000000000000010000000001; // D (0x0000000000000401) 
//    12'ha54 : errs =          63'b000000000000000000000000000000000000000000000000000100000000001; // D (0x0000000000000801) 
//    12'heda : errs =          63'b000000000000000000000000000000000000000000000000001000000000001; // D (0x0000000000001001) 
//    12'h7c6 : errs =          63'b000000000000000000000000000000000000000000000000010000000000001; // D (0x0000000000002001) 
//    12'h0c7 : errs =          63'b000000000000000000000000000000000000000000000000100000000000001; // D (0x0000000000004001) 
//    12'hec5 : errs =          63'b000000000000000000000000000000000000000000000001000000000000001; // D (0x0000000000008001) 
//    12'h7f8 : errs =          63'b000000000000000000000000000000000000000000000010000000000000001; // D (0x0000000000010001) 
//    12'h0bb : errs =          63'b000000000000000000000000000000000000000000000100000000000000001; // D (0x0000000000020001) 
//    12'he3d : errs =          63'b000000000000000000000000000000000000000000001000000000000000001; // D (0x0000000000040001) 
//    12'h608 : errs =          63'b000000000000000000000000000000000000000000010000000000000000001; // D (0x0000000000080001) 
//    12'h35b : errs =          63'b000000000000000000000000000000000000000000100000000000000000001; // D (0x0000000000100001) 
//    12'h9fd : errs =          63'b000000000000000000000000000000000000000001000000000000000000001; // D (0x0000000000200001) 
//    12'h988 : errs =          63'b000000000000000000000000000000000000000010000000000000000000001; // D (0x0000000000400001) 
//    12'h962 : errs =          63'b000000000000000000000000000000000000000100000000000000000000001; // D (0x0000000000800001) 
//    12'h8b6 : errs =          63'b000000000000000000000000000000000000001000000000000000000000001; // D (0x0000000001000001) 
//    12'hb1e : errs =          63'b000000000000000000000000000000000000010000000000000000000000001; // D (0x0000000002000001) 
//    12'hc4e : errs =          63'b000000000000000000000000000000000000100000000000000000000000001; // D (0x0000000004000001) 
//    12'h2ee : errs =          63'b000000000000000000000000000000000001000000000000000000000000001; // D (0x0000000008000001) 
//    12'ha97 : errs =          63'b000000000000000000000000000000000010000000000000000000000000001; // D (0x0000000010000001) 
//    12'hf5c : errs =          63'b000000000000000000000000000000000100000000000000000000000000001; // D (0x0000000020000001) 
//    12'h4ca : errs =          63'b000000000000000000000000000000001000000000000000000000000000001; // D (0x0000000040000001) 
//    12'h6df : errs =          63'b000000000000000000000000000000010000000000000000000000000000001; // D (0x0000000080000001) 
//    12'h2f5 : errs =          63'b000000000000000000000000000000100000000000000000000000000000001; // D (0x0000000100000001) 
//    12'haa1 : errs =          63'b000000000000000000000000000001000000000000000000000000000000001; // D (0x0000000200000001) 
//    12'hf30 : errs =          63'b000000000000000000000000000010000000000000000000000000000000001; // D (0x0000000400000001) 
//    12'h412 : errs =          63'b000000000000000000000000000100000000000000000000000000000000001; // D (0x0000000800000001) 
//    12'h76f : errs =          63'b000000000000000000000000001000000000000000000000000000000000001; // D (0x0000001000000001) 
//    12'h195 : errs =          63'b000000000000000000000000010000000000000000000000000000000000001; // D (0x0000002000000001) 
//    12'hc61 : errs =          63'b000000000000000000000000100000000000000000000000000000000000001; // D (0x0000004000000001) 
//    12'h2b0 : errs =          63'b000000000000000000000001000000000000000000000000000000000000001; // D (0x0000008000000001) 
//    12'ha2b : errs =          63'b000000000000000000000010000000000000000000000000000000000000001; // D (0x0000010000000001) 
//    12'he24 : errs =          63'b000000000000000000000100000000000000000000000000000000000000001; // D (0x0000020000000001) 
//    12'h63a : errs =          63'b000000000000000000001000000000000000000000000000000000000000001; // D (0x0000040000000001) 
//    12'h33f : errs =          63'b000000000000000000010000000000000000000000000000000000000000001; // D (0x0000080000000001) 
//    12'h935 : errs =          63'b000000000000000000100000000000000000000000000000000000000000001; // D (0x0000100000000001) 
//    12'h818 : errs =          63'b000000000000000001000000000000000000000000000000000000000000001; // D (0x0000200000000001) 
//    12'ha42 : errs =          63'b000000000000000010000000000000000000000000000000000000000000001; // D (0x0000400000000001) 
//    12'hef6 : errs =          63'b000000000000000100000000000000000000000000000000000000000000001; // D (0x0000800000000001) 
//    12'h79e : errs =          63'b000000000000001000000000000000000000000000000000000000000000001; // D (0x0001000000000001) 
//    12'h077 : errs =          63'b000000000000010000000000000000000000000000000000000000000000001; // D (0x0002000000000001) 
//    12'hfa5 : errs =          63'b000000000000100000000000000000000000000000000000000000000000001; // D (0x0004000000000001) 
//    12'h538 : errs =          63'b000000000001000000000000000000000000000000000000000000000000001; // D (0x0008000000000001) 
//    12'h53b : errs =          63'b000000000010000000000000000000000000000000000000000000000000001; // D (0x0010000000000001) 
//    12'h53d : errs =          63'b000000000100000000000000000000000000000000000000000000000000001; // D (0x0020000000000001) 
//    12'h531 : errs =          63'b000000001000000000000000000000000000000000000000000000000000001; // D (0x0040000000000001) 
//    12'h529 : errs =          63'b000000010000000000000000000000000000000000000000000000000000001; // D (0x0080000000000001) 
//    12'h519 : errs =          63'b000000100000000000000000000000000000000000000000000000000000001; // D (0x0100000000000001) 
//    12'h579 : errs =          63'b000001000000000000000000000000000000000000000000000000000000001; // D (0x0200000000000001) 
//    12'h5b9 : errs =          63'b000010000000000000000000000000000000000000000000000000000000001; // D (0x0400000000000001) 
//    12'h439 : errs =          63'b000100000000000000000000000000000000000000000000000000000000001; // D (0x0800000000000001) 
//    12'h739 : errs =          63'b001000000000000000000000000000000000000000000000000000000000001; // D (0x1000000000000001) 
//    12'h139 : errs =          63'b010000000000000000000000000000000000000000000000000000000000001; // D (0x2000000000000001) 
//    12'hd39 : errs =          63'b100000000000000000000000000000000000000000000000000000000000001; // D (0x4000000000000001) 
    12'hf4b : errs =          63'b000000000000000000000000000000000000000000000000000000000000011; // D (0x0000000000000003) 
    12'ha72 : errs =          63'b000000000000000000000000000000000000000000000000000000000000010; // S (0x0000000000000002) 
//    12'hbaf : errs =          63'b000000000000000000000000000000000000000000000000000000000000110; // D (0x0000000000000006) 
//    12'h9c8 : errs =          63'b000000000000000000000000000000000000000000000000000000000001010; // D (0x000000000000000a) 
//    12'hd06 : errs =          63'b000000000000000000000000000000000000000000000000000000000010010; // D (0x0000000000000012) 
//    12'h49a : errs =          63'b000000000000000000000000000000000000000000000000000000000100010; // D (0x0000000000000022) 
//    12'h29b : errs =          63'b000000000000000000000000000000000000000000000000000000001000010; // D (0x0000000000000042) 
//    12'he99 : errs =          63'b000000000000000000000000000000000000000000000000000000010000010; // D (0x0000000000000082) 
//    12'h3a4 : errs =          63'b000000000000000000000000000000000000000000000000000000100000010; // D (0x0000000000000102) 
//    12'hce7 : errs =          63'b000000000000000000000000000000000000000000000000000001000000010; // D (0x0000000000000202) 
//    12'h758 : errs =          63'b000000000000000000000000000000000000000000000000000010000000010; // D (0x0000000000000402) 
//    12'h51f : errs =          63'b000000000000000000000000000000000000000000000000000100000000010; // D (0x0000000000000802) 
//    12'h191 : errs =          63'b000000000000000000000000000000000000000000000000001000000000010; // D (0x0000000000001002) 
//    12'h88d : errs =          63'b000000000000000000000000000000000000000000000000010000000000010; // D (0x0000000000002002) 
//    12'hf8c : errs =          63'b000000000000000000000000000000000000000000000000100000000000010; // D (0x0000000000004002) 
//    12'h18e : errs =          63'b000000000000000000000000000000000000000000000001000000000000010; // D (0x0000000000008002) 
//    12'h8b3 : errs =          63'b000000000000000000000000000000000000000000000010000000000000010; // D (0x0000000000010002) 
//    12'hff0 : errs =          63'b000000000000000000000000000000000000000000000100000000000000010; // D (0x0000000000020002) 
//    12'h176 : errs =          63'b000000000000000000000000000000000000000000001000000000000000010; // D (0x0000000000040002) 
//    12'h943 : errs =          63'b000000000000000000000000000000000000000000010000000000000000010; // D (0x0000000000080002) 
//    12'hc10 : errs =          63'b000000000000000000000000000000000000000000100000000000000000010; // D (0x0000000000100002) 
//    12'h6b6 : errs =          63'b000000000000000000000000000000000000000001000000000000000000010; // D (0x0000000000200002) 
//    12'h6c3 : errs =          63'b000000000000000000000000000000000000000010000000000000000000010; // D (0x0000000000400002) 
//    12'h629 : errs =          63'b000000000000000000000000000000000000000100000000000000000000010; // D (0x0000000000800002) 
//    12'h7fd : errs =          63'b000000000000000000000000000000000000001000000000000000000000010; // D (0x0000000001000002) 
//    12'h455 : errs =          63'b000000000000000000000000000000000000010000000000000000000000010; // D (0x0000000002000002) 
//    12'h305 : errs =          63'b000000000000000000000000000000000000100000000000000000000000010; // D (0x0000000004000002) 
//    12'hda5 : errs =          63'b000000000000000000000000000000000001000000000000000000000000010; // D (0x0000000008000002) 
//    12'h5dc : errs =          63'b000000000000000000000000000000000010000000000000000000000000010; // D (0x0000000010000002) 
//    12'h017 : errs =          63'b000000000000000000000000000000000100000000000000000000000000010; // D (0x0000000020000002) 
//    12'hb81 : errs =          63'b000000000000000000000000000000001000000000000000000000000000010; // D (0x0000000040000002) 
//    12'h994 : errs =          63'b000000000000000000000000000000010000000000000000000000000000010; // D (0x0000000080000002) 
//    12'hdbe : errs =          63'b000000000000000000000000000000100000000000000000000000000000010; // D (0x0000000100000002) 
//    12'h5ea : errs =          63'b000000000000000000000000000001000000000000000000000000000000010; // D (0x0000000200000002) 
//    12'h07b : errs =          63'b000000000000000000000000000010000000000000000000000000000000010; // D (0x0000000400000002) 
//    12'hb59 : errs =          63'b000000000000000000000000000100000000000000000000000000000000010; // D (0x0000000800000002) 
//    12'h824 : errs =          63'b000000000000000000000000001000000000000000000000000000000000010; // D (0x0000001000000002) 
//    12'hede : errs =          63'b000000000000000000000000010000000000000000000000000000000000010; // D (0x0000002000000002) 
//    12'h32a : errs =          63'b000000000000000000000000100000000000000000000000000000000000010; // D (0x0000004000000002) 
//    12'hdfb : errs =          63'b000000000000000000000001000000000000000000000000000000000000010; // D (0x0000008000000002) 
//    12'h560 : errs =          63'b000000000000000000000010000000000000000000000000000000000000010; // D (0x0000010000000002) 
//    12'h16f : errs =          63'b000000000000000000000100000000000000000000000000000000000000010; // D (0x0000020000000002) 
//    12'h971 : errs =          63'b000000000000000000001000000000000000000000000000000000000000010; // D (0x0000040000000002) 
//    12'hc74 : errs =          63'b000000000000000000010000000000000000000000000000000000000000010; // D (0x0000080000000002) 
//    12'h67e : errs =          63'b000000000000000000100000000000000000000000000000000000000000010; // D (0x0000100000000002) 
//    12'h753 : errs =          63'b000000000000000001000000000000000000000000000000000000000000010; // D (0x0000200000000002) 
//    12'h509 : errs =          63'b000000000000000010000000000000000000000000000000000000000000010; // D (0x0000400000000002) 
//    12'h1bd : errs =          63'b000000000000000100000000000000000000000000000000000000000000010; // D (0x0000800000000002) 
//    12'h8d5 : errs =          63'b000000000000001000000000000000000000000000000000000000000000010; // D (0x0001000000000002) 
//    12'hf3c : errs =          63'b000000000000010000000000000000000000000000000000000000000000010; // D (0x0002000000000002) 
//    12'h0ee : errs =          63'b000000000000100000000000000000000000000000000000000000000000010; // D (0x0004000000000002) 
//    12'ha73 : errs =          63'b000000000001000000000000000000000000000000000000000000000000010; // D (0x0008000000000002) 
//    12'ha70 : errs =          63'b000000000010000000000000000000000000000000000000000000000000010; // D (0x0010000000000002) 
//    12'ha76 : errs =          63'b000000000100000000000000000000000000000000000000000000000000010; // D (0x0020000000000002) 
//    12'ha7a : errs =          63'b000000001000000000000000000000000000000000000000000000000000010; // D (0x0040000000000002) 
//    12'ha62 : errs =          63'b000000010000000000000000000000000000000000000000000000000000010; // D (0x0080000000000002) 
//    12'ha52 : errs =          63'b000000100000000000000000000000000000000000000000000000000000010; // D (0x0100000000000002) 
//    12'ha32 : errs =          63'b000001000000000000000000000000000000000000000000000000000000010; // D (0x0200000000000002) 
//    12'haf2 : errs =          63'b000010000000000000000000000000000000000000000000000000000000010; // D (0x0400000000000002) 
//    12'hb72 : errs =          63'b000100000000000000000000000000000000000000000000000000000000010; // D (0x0800000000000002) 
//    12'h872 : errs =          63'b001000000000000000000000000000000000000000000000000000000000010; // D (0x1000000000000002) 
//    12'he72 : errs =          63'b010000000000000000000000000000000000000000000000000000000000010; // D (0x2000000000000002) 
//    12'h272 : errs =          63'b100000000000000000000000000000000000000000000000000000000000010; // D (0x4000000000000002) 
    12'h4e4 : errs =          63'b000000000000000000000000000000000000000000000000000000000000101; // D (0x0000000000000005) 
    12'hbaf : errs =          63'b000000000000000000000000000000000000000000000000000000000000110; // D (0x0000000000000006) 
    12'h1dd : errs =          63'b000000000000000000000000000000000000000000000000000000000000100; // S (0x0000000000000004) 
//    12'h267 : errs =          63'b000000000000000000000000000000000000000000000000000000000001100; // D (0x000000000000000c) 
//    12'h6a9 : errs =          63'b000000000000000000000000000000000000000000000000000000000010100; // D (0x0000000000000014) 
//    12'hf35 : errs =          63'b000000000000000000000000000000000000000000000000000000000100100; // D (0x0000000000000024) 
//    12'h934 : errs =          63'b000000000000000000000000000000000000000000000000000000001000100; // D (0x0000000000000044) 
//    12'h536 : errs =          63'b000000000000000000000000000000000000000000000000000000010000100; // D (0x0000000000000084) 
//    12'h80b : errs =          63'b000000000000000000000000000000000000000000000000000000100000100; // D (0x0000000000000104) 
//    12'h748 : errs =          63'b000000000000000000000000000000000000000000000000000001000000100; // D (0x0000000000000204) 
//    12'hcf7 : errs =          63'b000000000000000000000000000000000000000000000000000010000000100; // D (0x0000000000000404) 
//    12'heb0 : errs =          63'b000000000000000000000000000000000000000000000000000100000000100; // D (0x0000000000000804) 
//    12'ha3e : errs =          63'b000000000000000000000000000000000000000000000000001000000000100; // D (0x0000000000001004) 
//    12'h322 : errs =          63'b000000000000000000000000000000000000000000000000010000000000100; // D (0x0000000000002004) 
//    12'h423 : errs =          63'b000000000000000000000000000000000000000000000000100000000000100; // D (0x0000000000004004) 
//    12'ha21 : errs =          63'b000000000000000000000000000000000000000000000001000000000000100; // D (0x0000000000008004) 
//    12'h31c : errs =          63'b000000000000000000000000000000000000000000000010000000000000100; // D (0x0000000000010004) 
//    12'h45f : errs =          63'b000000000000000000000000000000000000000000000100000000000000100; // D (0x0000000000020004) 
//    12'had9 : errs =          63'b000000000000000000000000000000000000000000001000000000000000100; // D (0x0000000000040004) 
//    12'h2ec : errs =          63'b000000000000000000000000000000000000000000010000000000000000100; // D (0x0000000000080004) 
//    12'h7bf : errs =          63'b000000000000000000000000000000000000000000100000000000000000100; // D (0x0000000000100004) 
//    12'hd19 : errs =          63'b000000000000000000000000000000000000000001000000000000000000100; // D (0x0000000000200004) 
//    12'hd6c : errs =          63'b000000000000000000000000000000000000000010000000000000000000100; // D (0x0000000000400004) 
//    12'hd86 : errs =          63'b000000000000000000000000000000000000000100000000000000000000100; // D (0x0000000000800004) 
//    12'hc52 : errs =          63'b000000000000000000000000000000000000001000000000000000000000100; // D (0x0000000001000004) 
//    12'hffa : errs =          63'b000000000000000000000000000000000000010000000000000000000000100; // D (0x0000000002000004) 
//    12'h8aa : errs =          63'b000000000000000000000000000000000000100000000000000000000000100; // D (0x0000000004000004) 
//    12'h60a : errs =          63'b000000000000000000000000000000000001000000000000000000000000100; // D (0x0000000008000004) 
//    12'he73 : errs =          63'b000000000000000000000000000000000010000000000000000000000000100; // D (0x0000000010000004) 
//    12'hbb8 : errs =          63'b000000000000000000000000000000000100000000000000000000000000100; // D (0x0000000020000004) 
//    12'h02e : errs =          63'b000000000000000000000000000000001000000000000000000000000000100; // D (0x0000000040000004) 
//    12'h23b : errs =          63'b000000000000000000000000000000010000000000000000000000000000100; // D (0x0000000080000004) 
//    12'h611 : errs =          63'b000000000000000000000000000000100000000000000000000000000000100; // D (0x0000000100000004) 
//    12'he45 : errs =          63'b000000000000000000000000000001000000000000000000000000000000100; // D (0x0000000200000004) 
//    12'hbd4 : errs =          63'b000000000000000000000000000010000000000000000000000000000000100; // D (0x0000000400000004) 
//    12'h0f6 : errs =          63'b000000000000000000000000000100000000000000000000000000000000100; // D (0x0000000800000004) 
//    12'h38b : errs =          63'b000000000000000000000000001000000000000000000000000000000000100; // D (0x0000001000000004) 
//    12'h571 : errs =          63'b000000000000000000000000010000000000000000000000000000000000100; // D (0x0000002000000004) 
//    12'h885 : errs =          63'b000000000000000000000000100000000000000000000000000000000000100; // D (0x0000004000000004) 
//    12'h654 : errs =          63'b000000000000000000000001000000000000000000000000000000000000100; // D (0x0000008000000004) 
//    12'hecf : errs =          63'b000000000000000000000010000000000000000000000000000000000000100; // D (0x0000010000000004) 
//    12'hac0 : errs =          63'b000000000000000000000100000000000000000000000000000000000000100; // D (0x0000020000000004) 
//    12'h2de : errs =          63'b000000000000000000001000000000000000000000000000000000000000100; // D (0x0000040000000004) 
//    12'h7db : errs =          63'b000000000000000000010000000000000000000000000000000000000000100; // D (0x0000080000000004) 
//    12'hdd1 : errs =          63'b000000000000000000100000000000000000000000000000000000000000100; // D (0x0000100000000004) 
//    12'hcfc : errs =          63'b000000000000000001000000000000000000000000000000000000000000100; // D (0x0000200000000004) 
//    12'hea6 : errs =          63'b000000000000000010000000000000000000000000000000000000000000100; // D (0x0000400000000004) 
//    12'ha12 : errs =          63'b000000000000000100000000000000000000000000000000000000000000100; // D (0x0000800000000004) 
//    12'h37a : errs =          63'b000000000000001000000000000000000000000000000000000000000000100; // D (0x0001000000000004) 
//    12'h493 : errs =          63'b000000000000010000000000000000000000000000000000000000000000100; // D (0x0002000000000004) 
//    12'hb41 : errs =          63'b000000000000100000000000000000000000000000000000000000000000100; // D (0x0004000000000004) 
//    12'h1dc : errs =          63'b000000000001000000000000000000000000000000000000000000000000100; // D (0x0008000000000004) 
//    12'h1df : errs =          63'b000000000010000000000000000000000000000000000000000000000000100; // D (0x0010000000000004) 
//    12'h1d9 : errs =          63'b000000000100000000000000000000000000000000000000000000000000100; // D (0x0020000000000004) 
//    12'h1d5 : errs =          63'b000000001000000000000000000000000000000000000000000000000000100; // D (0x0040000000000004) 
//    12'h1cd : errs =          63'b000000010000000000000000000000000000000000000000000000000000100; // D (0x0080000000000004) 
//    12'h1fd : errs =          63'b000000100000000000000000000000000000000000000000000000000000100; // D (0x0100000000000004) 
//    12'h19d : errs =          63'b000001000000000000000000000000000000000000000000000000000000100; // D (0x0200000000000004) 
//    12'h15d : errs =          63'b000010000000000000000000000000000000000000000000000000000000100; // D (0x0400000000000004) 
//    12'h0dd : errs =          63'b000100000000000000000000000000000000000000000000000000000000100; // D (0x0800000000000004) 
//    12'h3dd : errs =          63'b001000000000000000000000000000000000000000000000000000000000100; // D (0x1000000000000004) 
//    12'h5dd : errs =          63'b010000000000000000000000000000000000000000000000000000000000100; // D (0x2000000000000004) 
//    12'h9dd : errs =          63'b100000000000000000000000000000000000000000000000000000000000100; // D (0x4000000000000004) 
    12'h683 : errs =          63'b000000000000000000000000000000000000000000000000000000000001001; // D (0x0000000000000009) 
    12'h9c8 : errs =          63'b000000000000000000000000000000000000000000000000000000000001010; // D (0x000000000000000a) 
    12'h267 : errs =          63'b000000000000000000000000000000000000000000000000000000000001100; // D (0x000000000000000c) 
    12'h3ba : errs =          63'b000000000000000000000000000000000000000000000000000000000001000; // S (0x0000000000000008) 
//    12'h4ce : errs =          63'b000000000000000000000000000000000000000000000000000000000011000; // D (0x0000000000000018) 
//    12'hd52 : errs =          63'b000000000000000000000000000000000000000000000000000000000101000; // D (0x0000000000000028) 
//    12'hb53 : errs =          63'b000000000000000000000000000000000000000000000000000000001001000; // D (0x0000000000000048) 
//    12'h751 : errs =          63'b000000000000000000000000000000000000000000000000000000010001000; // D (0x0000000000000088) 
//    12'ha6c : errs =          63'b000000000000000000000000000000000000000000000000000000100001000; // D (0x0000000000000108) 
//    12'h52f : errs =          63'b000000000000000000000000000000000000000000000000000001000001000; // D (0x0000000000000208) 
//    12'he90 : errs =          63'b000000000000000000000000000000000000000000000000000010000001000; // D (0x0000000000000408) 
//    12'hcd7 : errs =          63'b000000000000000000000000000000000000000000000000000100000001000; // D (0x0000000000000808) 
//    12'h859 : errs =          63'b000000000000000000000000000000000000000000000000001000000001000; // D (0x0000000000001008) 
//    12'h145 : errs =          63'b000000000000000000000000000000000000000000000000010000000001000; // D (0x0000000000002008) 
//    12'h644 : errs =          63'b000000000000000000000000000000000000000000000000100000000001000; // D (0x0000000000004008) 
//    12'h846 : errs =          63'b000000000000000000000000000000000000000000000001000000000001000; // D (0x0000000000008008) 
//    12'h17b : errs =          63'b000000000000000000000000000000000000000000000010000000000001000; // D (0x0000000000010008) 
//    12'h638 : errs =          63'b000000000000000000000000000000000000000000000100000000000001000; // D (0x0000000000020008) 
//    12'h8be : errs =          63'b000000000000000000000000000000000000000000001000000000000001000; // D (0x0000000000040008) 
//    12'h08b : errs =          63'b000000000000000000000000000000000000000000010000000000000001000; // D (0x0000000000080008) 
//    12'h5d8 : errs =          63'b000000000000000000000000000000000000000000100000000000000001000; // D (0x0000000000100008) 
//    12'hf7e : errs =          63'b000000000000000000000000000000000000000001000000000000000001000; // D (0x0000000000200008) 
//    12'hf0b : errs =          63'b000000000000000000000000000000000000000010000000000000000001000; // D (0x0000000000400008) 
//    12'hfe1 : errs =          63'b000000000000000000000000000000000000000100000000000000000001000; // D (0x0000000000800008) 
//    12'he35 : errs =          63'b000000000000000000000000000000000000001000000000000000000001000; // D (0x0000000001000008) 
//    12'hd9d : errs =          63'b000000000000000000000000000000000000010000000000000000000001000; // D (0x0000000002000008) 
//    12'hacd : errs =          63'b000000000000000000000000000000000000100000000000000000000001000; // D (0x0000000004000008) 
//    12'h46d : errs =          63'b000000000000000000000000000000000001000000000000000000000001000; // D (0x0000000008000008) 
//    12'hc14 : errs =          63'b000000000000000000000000000000000010000000000000000000000001000; // D (0x0000000010000008) 
//    12'h9df : errs =          63'b000000000000000000000000000000000100000000000000000000000001000; // D (0x0000000020000008) 
//    12'h249 : errs =          63'b000000000000000000000000000000001000000000000000000000000001000; // D (0x0000000040000008) 
//    12'h05c : errs =          63'b000000000000000000000000000000010000000000000000000000000001000; // D (0x0000000080000008) 
//    12'h476 : errs =          63'b000000000000000000000000000000100000000000000000000000000001000; // D (0x0000000100000008) 
//    12'hc22 : errs =          63'b000000000000000000000000000001000000000000000000000000000001000; // D (0x0000000200000008) 
//    12'h9b3 : errs =          63'b000000000000000000000000000010000000000000000000000000000001000; // D (0x0000000400000008) 
//    12'h291 : errs =          63'b000000000000000000000000000100000000000000000000000000000001000; // D (0x0000000800000008) 
//    12'h1ec : errs =          63'b000000000000000000000000001000000000000000000000000000000001000; // D (0x0000001000000008) 
//    12'h716 : errs =          63'b000000000000000000000000010000000000000000000000000000000001000; // D (0x0000002000000008) 
//    12'hae2 : errs =          63'b000000000000000000000000100000000000000000000000000000000001000; // D (0x0000004000000008) 
//    12'h433 : errs =          63'b000000000000000000000001000000000000000000000000000000000001000; // D (0x0000008000000008) 
//    12'hca8 : errs =          63'b000000000000000000000010000000000000000000000000000000000001000; // D (0x0000010000000008) 
//    12'h8a7 : errs =          63'b000000000000000000000100000000000000000000000000000000000001000; // D (0x0000020000000008) 
//    12'h0b9 : errs =          63'b000000000000000000001000000000000000000000000000000000000001000; // D (0x0000040000000008) 
//    12'h5bc : errs =          63'b000000000000000000010000000000000000000000000000000000000001000; // D (0x0000080000000008) 
//    12'hfb6 : errs =          63'b000000000000000000100000000000000000000000000000000000000001000; // D (0x0000100000000008) 
//    12'he9b : errs =          63'b000000000000000001000000000000000000000000000000000000000001000; // D (0x0000200000000008) 
//    12'hcc1 : errs =          63'b000000000000000010000000000000000000000000000000000000000001000; // D (0x0000400000000008) 
//    12'h875 : errs =          63'b000000000000000100000000000000000000000000000000000000000001000; // D (0x0000800000000008) 
//    12'h11d : errs =          63'b000000000000001000000000000000000000000000000000000000000001000; // D (0x0001000000000008) 
//    12'h6f4 : errs =          63'b000000000000010000000000000000000000000000000000000000000001000; // D (0x0002000000000008) 
//    12'h926 : errs =          63'b000000000000100000000000000000000000000000000000000000000001000; // D (0x0004000000000008) 
//    12'h3bb : errs =          63'b000000000001000000000000000000000000000000000000000000000001000; // D (0x0008000000000008) 
//    12'h3b8 : errs =          63'b000000000010000000000000000000000000000000000000000000000001000; // D (0x0010000000000008) 
//    12'h3be : errs =          63'b000000000100000000000000000000000000000000000000000000000001000; // D (0x0020000000000008) 
//    12'h3b2 : errs =          63'b000000001000000000000000000000000000000000000000000000000001000; // D (0x0040000000000008) 
//    12'h3aa : errs =          63'b000000010000000000000000000000000000000000000000000000000001000; // D (0x0080000000000008) 
//    12'h39a : errs =          63'b000000100000000000000000000000000000000000000000000000000001000; // D (0x0100000000000008) 
//    12'h3fa : errs =          63'b000001000000000000000000000000000000000000000000000000000001000; // D (0x0200000000000008) 
//    12'h33a : errs =          63'b000010000000000000000000000000000000000000000000000000000001000; // D (0x0400000000000008) 
//    12'h2ba : errs =          63'b000100000000000000000000000000000000000000000000000000000001000; // D (0x0800000000000008) 
//    12'h1ba : errs =          63'b001000000000000000000000000000000000000000000000000000000001000; // D (0x1000000000000008) 
//    12'h7ba : errs =          63'b010000000000000000000000000000000000000000000000000000000001000; // D (0x2000000000000008) 
//    12'hbba : errs =          63'b100000000000000000000000000000000000000000000000000000000001000; // D (0x4000000000000008) 
    12'h24d : errs =          63'b000000000000000000000000000000000000000000000000000000000010001; // D (0x0000000000000011) 
    12'hd06 : errs =          63'b000000000000000000000000000000000000000000000000000000000010010; // D (0x0000000000000012) 
    12'h6a9 : errs =          63'b000000000000000000000000000000000000000000000000000000000010100; // D (0x0000000000000014) 
    12'h4ce : errs =          63'b000000000000000000000000000000000000000000000000000000000011000; // D (0x0000000000000018) 
    12'h774 : errs =          63'b000000000000000000000000000000000000000000000000000000000010000; // S (0x0000000000000010) 
//    12'h99c : errs =          63'b000000000000000000000000000000000000000000000000000000000110000; // D (0x0000000000000030) 
//    12'hf9d : errs =          63'b000000000000000000000000000000000000000000000000000000001010000; // D (0x0000000000000050) 
//    12'h39f : errs =          63'b000000000000000000000000000000000000000000000000000000010010000; // D (0x0000000000000090) 
//    12'hea2 : errs =          63'b000000000000000000000000000000000000000000000000000000100010000; // D (0x0000000000000110) 
//    12'h1e1 : errs =          63'b000000000000000000000000000000000000000000000000000001000010000; // D (0x0000000000000210) 
//    12'ha5e : errs =          63'b000000000000000000000000000000000000000000000000000010000010000; // D (0x0000000000000410) 
//    12'h819 : errs =          63'b000000000000000000000000000000000000000000000000000100000010000; // D (0x0000000000000810) 
//    12'hc97 : errs =          63'b000000000000000000000000000000000000000000000000001000000010000; // D (0x0000000000001010) 
//    12'h58b : errs =          63'b000000000000000000000000000000000000000000000000010000000010000; // D (0x0000000000002010) 
//    12'h28a : errs =          63'b000000000000000000000000000000000000000000000000100000000010000; // D (0x0000000000004010) 
//    12'hc88 : errs =          63'b000000000000000000000000000000000000000000000001000000000010000; // D (0x0000000000008010) 
//    12'h5b5 : errs =          63'b000000000000000000000000000000000000000000000010000000000010000; // D (0x0000000000010010) 
//    12'h2f6 : errs =          63'b000000000000000000000000000000000000000000000100000000000010000; // D (0x0000000000020010) 
//    12'hc70 : errs =          63'b000000000000000000000000000000000000000000001000000000000010000; // D (0x0000000000040010) 
//    12'h445 : errs =          63'b000000000000000000000000000000000000000000010000000000000010000; // D (0x0000000000080010) 
//    12'h116 : errs =          63'b000000000000000000000000000000000000000000100000000000000010000; // D (0x0000000000100010) 
//    12'hbb0 : errs =          63'b000000000000000000000000000000000000000001000000000000000010000; // D (0x0000000000200010) 
//    12'hbc5 : errs =          63'b000000000000000000000000000000000000000010000000000000000010000; // D (0x0000000000400010) 
//    12'hb2f : errs =          63'b000000000000000000000000000000000000000100000000000000000010000; // D (0x0000000000800010) 
//    12'hafb : errs =          63'b000000000000000000000000000000000000001000000000000000000010000; // D (0x0000000001000010) 
//    12'h953 : errs =          63'b000000000000000000000000000000000000010000000000000000000010000; // D (0x0000000002000010) 
//    12'he03 : errs =          63'b000000000000000000000000000000000000100000000000000000000010000; // D (0x0000000004000010) 
//    12'h0a3 : errs =          63'b000000000000000000000000000000000001000000000000000000000010000; // D (0x0000000008000010) 
//    12'h8da : errs =          63'b000000000000000000000000000000000010000000000000000000000010000; // D (0x0000000010000010) 
//    12'hd11 : errs =          63'b000000000000000000000000000000000100000000000000000000000010000; // D (0x0000000020000010) 
//    12'h687 : errs =          63'b000000000000000000000000000000001000000000000000000000000010000; // D (0x0000000040000010) 
//    12'h492 : errs =          63'b000000000000000000000000000000010000000000000000000000000010000; // D (0x0000000080000010) 
//    12'h0b8 : errs =          63'b000000000000000000000000000000100000000000000000000000000010000; // D (0x0000000100000010) 
//    12'h8ec : errs =          63'b000000000000000000000000000001000000000000000000000000000010000; // D (0x0000000200000010) 
//    12'hd7d : errs =          63'b000000000000000000000000000010000000000000000000000000000010000; // D (0x0000000400000010) 
//    12'h65f : errs =          63'b000000000000000000000000000100000000000000000000000000000010000; // D (0x0000000800000010) 
//    12'h522 : errs =          63'b000000000000000000000000001000000000000000000000000000000010000; // D (0x0000001000000010) 
//    12'h3d8 : errs =          63'b000000000000000000000000010000000000000000000000000000000010000; // D (0x0000002000000010) 
//    12'he2c : errs =          63'b000000000000000000000000100000000000000000000000000000000010000; // D (0x0000004000000010) 
//    12'h0fd : errs =          63'b000000000000000000000001000000000000000000000000000000000010000; // D (0x0000008000000010) 
//    12'h866 : errs =          63'b000000000000000000000010000000000000000000000000000000000010000; // D (0x0000010000000010) 
//    12'hc69 : errs =          63'b000000000000000000000100000000000000000000000000000000000010000; // D (0x0000020000000010) 
//    12'h477 : errs =          63'b000000000000000000001000000000000000000000000000000000000010000; // D (0x0000040000000010) 
//    12'h172 : errs =          63'b000000000000000000010000000000000000000000000000000000000010000; // D (0x0000080000000010) 
//    12'hb78 : errs =          63'b000000000000000000100000000000000000000000000000000000000010000; // D (0x0000100000000010) 
//    12'ha55 : errs =          63'b000000000000000001000000000000000000000000000000000000000010000; // D (0x0000200000000010) 
//    12'h80f : errs =          63'b000000000000000010000000000000000000000000000000000000000010000; // D (0x0000400000000010) 
//    12'hcbb : errs =          63'b000000000000000100000000000000000000000000000000000000000010000; // D (0x0000800000000010) 
//    12'h5d3 : errs =          63'b000000000000001000000000000000000000000000000000000000000010000; // D (0x0001000000000010) 
//    12'h23a : errs =          63'b000000000000010000000000000000000000000000000000000000000010000; // D (0x0002000000000010) 
//    12'hde8 : errs =          63'b000000000000100000000000000000000000000000000000000000000010000; // D (0x0004000000000010) 
//    12'h775 : errs =          63'b000000000001000000000000000000000000000000000000000000000010000; // D (0x0008000000000010) 
//    12'h776 : errs =          63'b000000000010000000000000000000000000000000000000000000000010000; // D (0x0010000000000010) 
//    12'h770 : errs =          63'b000000000100000000000000000000000000000000000000000000000010000; // D (0x0020000000000010) 
//    12'h77c : errs =          63'b000000001000000000000000000000000000000000000000000000000010000; // D (0x0040000000000010) 
//    12'h764 : errs =          63'b000000010000000000000000000000000000000000000000000000000010000; // D (0x0080000000000010) 
//    12'h754 : errs =          63'b000000100000000000000000000000000000000000000000000000000010000; // D (0x0100000000000010) 
//    12'h734 : errs =          63'b000001000000000000000000000000000000000000000000000000000010000; // D (0x0200000000000010) 
//    12'h7f4 : errs =          63'b000010000000000000000000000000000000000000000000000000000010000; // D (0x0400000000000010) 
//    12'h674 : errs =          63'b000100000000000000000000000000000000000000000000000000000010000; // D (0x0800000000000010) 
//    12'h574 : errs =          63'b001000000000000000000000000000000000000000000000000000000010000; // D (0x1000000000000010) 
//    12'h374 : errs =          63'b010000000000000000000000000000000000000000000000000000000010000; // D (0x2000000000000010) 
//    12'hf74 : errs =          63'b100000000000000000000000000000000000000000000000000000000010000; // D (0x4000000000000010) 
    12'hbd1 : errs =          63'b000000000000000000000000000000000000000000000000000000000100001; // D (0x0000000000000021) 
    12'h49a : errs =          63'b000000000000000000000000000000000000000000000000000000000100010; // D (0x0000000000000022) 
    12'hf35 : errs =          63'b000000000000000000000000000000000000000000000000000000000100100; // D (0x0000000000000024) 
    12'hd52 : errs =          63'b000000000000000000000000000000000000000000000000000000000101000; // D (0x0000000000000028) 
    12'h99c : errs =          63'b000000000000000000000000000000000000000000000000000000000110000; // D (0x0000000000000030) 
    12'hee8 : errs =          63'b000000000000000000000000000000000000000000000000000000000100000; // S (0x0000000000000020) 
//    12'h601 : errs =          63'b000000000000000000000000000000000000000000000000000000001100000; // D (0x0000000000000060) 
//    12'ha03 : errs =          63'b000000000000000000000000000000000000000000000000000000010100000; // D (0x00000000000000a0) 
//    12'h73e : errs =          63'b000000000000000000000000000000000000000000000000000000100100000; // D (0x0000000000000120) 
//    12'h87d : errs =          63'b000000000000000000000000000000000000000000000000000001000100000; // D (0x0000000000000220) 
//    12'h3c2 : errs =          63'b000000000000000000000000000000000000000000000000000010000100000; // D (0x0000000000000420) 
//    12'h185 : errs =          63'b000000000000000000000000000000000000000000000000000100000100000; // D (0x0000000000000820) 
//    12'h50b : errs =          63'b000000000000000000000000000000000000000000000000001000000100000; // D (0x0000000000001020) 
//    12'hc17 : errs =          63'b000000000000000000000000000000000000000000000000010000000100000; // D (0x0000000000002020) 
//    12'hb16 : errs =          63'b000000000000000000000000000000000000000000000000100000000100000; // D (0x0000000000004020) 
//    12'h514 : errs =          63'b000000000000000000000000000000000000000000000001000000000100000; // D (0x0000000000008020) 
//    12'hc29 : errs =          63'b000000000000000000000000000000000000000000000010000000000100000; // D (0x0000000000010020) 
//    12'hb6a : errs =          63'b000000000000000000000000000000000000000000000100000000000100000; // D (0x0000000000020020) 
//    12'h5ec : errs =          63'b000000000000000000000000000000000000000000001000000000000100000; // D (0x0000000000040020) 
//    12'hdd9 : errs =          63'b000000000000000000000000000000000000000000010000000000000100000; // D (0x0000000000080020) 
//    12'h88a : errs =          63'b000000000000000000000000000000000000000000100000000000000100000; // D (0x0000000000100020) 
//    12'h22c : errs =          63'b000000000000000000000000000000000000000001000000000000000100000; // D (0x0000000000200020) 
//    12'h259 : errs =          63'b000000000000000000000000000000000000000010000000000000000100000; // D (0x0000000000400020) 
//    12'h2b3 : errs =          63'b000000000000000000000000000000000000000100000000000000000100000; // D (0x0000000000800020) 
//    12'h367 : errs =          63'b000000000000000000000000000000000000001000000000000000000100000; // D (0x0000000001000020) 
//    12'h0cf : errs =          63'b000000000000000000000000000000000000010000000000000000000100000; // D (0x0000000002000020) 
//    12'h79f : errs =          63'b000000000000000000000000000000000000100000000000000000000100000; // D (0x0000000004000020) 
//    12'h93f : errs =          63'b000000000000000000000000000000000001000000000000000000000100000; // D (0x0000000008000020) 
//    12'h146 : errs =          63'b000000000000000000000000000000000010000000000000000000000100000; // D (0x0000000010000020) 
//    12'h48d : errs =          63'b000000000000000000000000000000000100000000000000000000000100000; // D (0x0000000020000020) 
//    12'hf1b : errs =          63'b000000000000000000000000000000001000000000000000000000000100000; // D (0x0000000040000020) 
//    12'hd0e : errs =          63'b000000000000000000000000000000010000000000000000000000000100000; // D (0x0000000080000020) 
//    12'h924 : errs =          63'b000000000000000000000000000000100000000000000000000000000100000; // D (0x0000000100000020) 
//    12'h170 : errs =          63'b000000000000000000000000000001000000000000000000000000000100000; // D (0x0000000200000020) 
//    12'h4e1 : errs =          63'b000000000000000000000000000010000000000000000000000000000100000; // D (0x0000000400000020) 
//    12'hfc3 : errs =          63'b000000000000000000000000000100000000000000000000000000000100000; // D (0x0000000800000020) 
//    12'hcbe : errs =          63'b000000000000000000000000001000000000000000000000000000000100000; // D (0x0000001000000020) 
//    12'ha44 : errs =          63'b000000000000000000000000010000000000000000000000000000000100000; // D (0x0000002000000020) 
//    12'h7b0 : errs =          63'b000000000000000000000000100000000000000000000000000000000100000; // D (0x0000004000000020) 
//    12'h961 : errs =          63'b000000000000000000000001000000000000000000000000000000000100000; // D (0x0000008000000020) 
//    12'h1fa : errs =          63'b000000000000000000000010000000000000000000000000000000000100000; // D (0x0000010000000020) 
//    12'h5f5 : errs =          63'b000000000000000000000100000000000000000000000000000000000100000; // D (0x0000020000000020) 
//    12'hdeb : errs =          63'b000000000000000000001000000000000000000000000000000000000100000; // D (0x0000040000000020) 
//    12'h8ee : errs =          63'b000000000000000000010000000000000000000000000000000000000100000; // D (0x0000080000000020) 
//    12'h2e4 : errs =          63'b000000000000000000100000000000000000000000000000000000000100000; // D (0x0000100000000020) 
//    12'h3c9 : errs =          63'b000000000000000001000000000000000000000000000000000000000100000; // D (0x0000200000000020) 
//    12'h193 : errs =          63'b000000000000000010000000000000000000000000000000000000000100000; // D (0x0000400000000020) 
//    12'h527 : errs =          63'b000000000000000100000000000000000000000000000000000000000100000; // D (0x0000800000000020) 
//    12'hc4f : errs =          63'b000000000000001000000000000000000000000000000000000000000100000; // D (0x0001000000000020) 
//    12'hba6 : errs =          63'b000000000000010000000000000000000000000000000000000000000100000; // D (0x0002000000000020) 
//    12'h474 : errs =          63'b000000000000100000000000000000000000000000000000000000000100000; // D (0x0004000000000020) 
//    12'hee9 : errs =          63'b000000000001000000000000000000000000000000000000000000000100000; // D (0x0008000000000020) 
//    12'heea : errs =          63'b000000000010000000000000000000000000000000000000000000000100000; // D (0x0010000000000020) 
//    12'heec : errs =          63'b000000000100000000000000000000000000000000000000000000000100000; // D (0x0020000000000020) 
//    12'hee0 : errs =          63'b000000001000000000000000000000000000000000000000000000000100000; // D (0x0040000000000020) 
//    12'hef8 : errs =          63'b000000010000000000000000000000000000000000000000000000000100000; // D (0x0080000000000020) 
//    12'hec8 : errs =          63'b000000100000000000000000000000000000000000000000000000000100000; // D (0x0100000000000020) 
//    12'hea8 : errs =          63'b000001000000000000000000000000000000000000000000000000000100000; // D (0x0200000000000020) 
//    12'he68 : errs =          63'b000010000000000000000000000000000000000000000000000000000100000; // D (0x0400000000000020) 
//    12'hfe8 : errs =          63'b000100000000000000000000000000000000000000000000000000000100000; // D (0x0800000000000020) 
//    12'hce8 : errs =          63'b001000000000000000000000000000000000000000000000000000000100000; // D (0x1000000000000020) 
//    12'hae8 : errs =          63'b010000000000000000000000000000000000000000000000000000000100000; // D (0x2000000000000020) 
//    12'h6e8 : errs =          63'b100000000000000000000000000000000000000000000000000000000100000; // D (0x4000000000000020) 
    12'hdd0 : errs =          63'b000000000000000000000000000000000000000000000000000000001000001; // D (0x0000000000000041) 
    12'h29b : errs =          63'b000000000000000000000000000000000000000000000000000000001000010; // D (0x0000000000000042) 
    12'h934 : errs =          63'b000000000000000000000000000000000000000000000000000000001000100; // D (0x0000000000000044) 
    12'hb53 : errs =          63'b000000000000000000000000000000000000000000000000000000001001000; // D (0x0000000000000048) 
    12'hf9d : errs =          63'b000000000000000000000000000000000000000000000000000000001010000; // D (0x0000000000000050) 
    12'h601 : errs =          63'b000000000000000000000000000000000000000000000000000000001100000; // D (0x0000000000000060) 
    12'h8e9 : errs =          63'b000000000000000000000000000000000000000000000000000000001000000; // S (0x0000000000000040) 
//    12'hc02 : errs =          63'b000000000000000000000000000000000000000000000000000000011000000; // D (0x00000000000000c0) 
//    12'h13f : errs =          63'b000000000000000000000000000000000000000000000000000000101000000; // D (0x0000000000000140) 
//    12'he7c : errs =          63'b000000000000000000000000000000000000000000000000000001001000000; // D (0x0000000000000240) 
//    12'h5c3 : errs =          63'b000000000000000000000000000000000000000000000000000010001000000; // D (0x0000000000000440) 
//    12'h784 : errs =          63'b000000000000000000000000000000000000000000000000000100001000000; // D (0x0000000000000840) 
//    12'h30a : errs =          63'b000000000000000000000000000000000000000000000000001000001000000; // D (0x0000000000001040) 
//    12'ha16 : errs =          63'b000000000000000000000000000000000000000000000000010000001000000; // D (0x0000000000002040) 
//    12'hd17 : errs =          63'b000000000000000000000000000000000000000000000000100000001000000; // D (0x0000000000004040) 
//    12'h315 : errs =          63'b000000000000000000000000000000000000000000000001000000001000000; // D (0x0000000000008040) 
//    12'ha28 : errs =          63'b000000000000000000000000000000000000000000000010000000001000000; // D (0x0000000000010040) 
//    12'hd6b : errs =          63'b000000000000000000000000000000000000000000000100000000001000000; // D (0x0000000000020040) 
//    12'h3ed : errs =          63'b000000000000000000000000000000000000000000001000000000001000000; // D (0x0000000000040040) 
//    12'hbd8 : errs =          63'b000000000000000000000000000000000000000000010000000000001000000; // D (0x0000000000080040) 
//    12'he8b : errs =          63'b000000000000000000000000000000000000000000100000000000001000000; // D (0x0000000000100040) 
//    12'h42d : errs =          63'b000000000000000000000000000000000000000001000000000000001000000; // D (0x0000000000200040) 
//    12'h458 : errs =          63'b000000000000000000000000000000000000000010000000000000001000000; // D (0x0000000000400040) 
//    12'h4b2 : errs =          63'b000000000000000000000000000000000000000100000000000000001000000; // D (0x0000000000800040) 
//    12'h566 : errs =          63'b000000000000000000000000000000000000001000000000000000001000000; // D (0x0000000001000040) 
//    12'h6ce : errs =          63'b000000000000000000000000000000000000010000000000000000001000000; // D (0x0000000002000040) 
//    12'h19e : errs =          63'b000000000000000000000000000000000000100000000000000000001000000; // D (0x0000000004000040) 
//    12'hf3e : errs =          63'b000000000000000000000000000000000001000000000000000000001000000; // D (0x0000000008000040) 
//    12'h747 : errs =          63'b000000000000000000000000000000000010000000000000000000001000000; // D (0x0000000010000040) 
//    12'h28c : errs =          63'b000000000000000000000000000000000100000000000000000000001000000; // D (0x0000000020000040) 
//    12'h91a : errs =          63'b000000000000000000000000000000001000000000000000000000001000000; // D (0x0000000040000040) 
//    12'hb0f : errs =          63'b000000000000000000000000000000010000000000000000000000001000000; // D (0x0000000080000040) 
//    12'hf25 : errs =          63'b000000000000000000000000000000100000000000000000000000001000000; // D (0x0000000100000040) 
//    12'h771 : errs =          63'b000000000000000000000000000001000000000000000000000000001000000; // D (0x0000000200000040) 
//    12'h2e0 : errs =          63'b000000000000000000000000000010000000000000000000000000001000000; // D (0x0000000400000040) 
//    12'h9c2 : errs =          63'b000000000000000000000000000100000000000000000000000000001000000; // D (0x0000000800000040) 
//    12'habf : errs =          63'b000000000000000000000000001000000000000000000000000000001000000; // D (0x0000001000000040) 
//    12'hc45 : errs =          63'b000000000000000000000000010000000000000000000000000000001000000; // D (0x0000002000000040) 
//    12'h1b1 : errs =          63'b000000000000000000000000100000000000000000000000000000001000000; // D (0x0000004000000040) 
//    12'hf60 : errs =          63'b000000000000000000000001000000000000000000000000000000001000000; // D (0x0000008000000040) 
//    12'h7fb : errs =          63'b000000000000000000000010000000000000000000000000000000001000000; // D (0x0000010000000040) 
//    12'h3f4 : errs =          63'b000000000000000000000100000000000000000000000000000000001000000; // D (0x0000020000000040) 
//    12'hbea : errs =          63'b000000000000000000001000000000000000000000000000000000001000000; // D (0x0000040000000040) 
//    12'heef : errs =          63'b000000000000000000010000000000000000000000000000000000001000000; // D (0x0000080000000040) 
//    12'h4e5 : errs =          63'b000000000000000000100000000000000000000000000000000000001000000; // D (0x0000100000000040) 
//    12'h5c8 : errs =          63'b000000000000000001000000000000000000000000000000000000001000000; // D (0x0000200000000040) 
//    12'h792 : errs =          63'b000000000000000010000000000000000000000000000000000000001000000; // D (0x0000400000000040) 
//    12'h326 : errs =          63'b000000000000000100000000000000000000000000000000000000001000000; // D (0x0000800000000040) 
//    12'ha4e : errs =          63'b000000000000001000000000000000000000000000000000000000001000000; // D (0x0001000000000040) 
//    12'hda7 : errs =          63'b000000000000010000000000000000000000000000000000000000001000000; // D (0x0002000000000040) 
//    12'h275 : errs =          63'b000000000000100000000000000000000000000000000000000000001000000; // D (0x0004000000000040) 
//    12'h8e8 : errs =          63'b000000000001000000000000000000000000000000000000000000001000000; // D (0x0008000000000040) 
//    12'h8eb : errs =          63'b000000000010000000000000000000000000000000000000000000001000000; // D (0x0010000000000040) 
//    12'h8ed : errs =          63'b000000000100000000000000000000000000000000000000000000001000000; // D (0x0020000000000040) 
//    12'h8e1 : errs =          63'b000000001000000000000000000000000000000000000000000000001000000; // D (0x0040000000000040) 
//    12'h8f9 : errs =          63'b000000010000000000000000000000000000000000000000000000001000000; // D (0x0080000000000040) 
//    12'h8c9 : errs =          63'b000000100000000000000000000000000000000000000000000000001000000; // D (0x0100000000000040) 
//    12'h8a9 : errs =          63'b000001000000000000000000000000000000000000000000000000001000000; // D (0x0200000000000040) 
//    12'h869 : errs =          63'b000010000000000000000000000000000000000000000000000000001000000; // D (0x0400000000000040) 
//    12'h9e9 : errs =          63'b000100000000000000000000000000000000000000000000000000001000000; // D (0x0800000000000040) 
//    12'hae9 : errs =          63'b001000000000000000000000000000000000000000000000000000001000000; // D (0x1000000000000040) 
//    12'hce9 : errs =          63'b010000000000000000000000000000000000000000000000000000001000000; // D (0x2000000000000040) 
//    12'h0e9 : errs =          63'b100000000000000000000000000000000000000000000000000000001000000; // D (0x4000000000000040) 
    12'h1d2 : errs =          63'b000000000000000000000000000000000000000000000000000000010000001; // D (0x0000000000000081) 
    12'he99 : errs =          63'b000000000000000000000000000000000000000000000000000000010000010; // D (0x0000000000000082) 
    12'h536 : errs =          63'b000000000000000000000000000000000000000000000000000000010000100; // D (0x0000000000000084) 
    12'h751 : errs =          63'b000000000000000000000000000000000000000000000000000000010001000; // D (0x0000000000000088) 
    12'h39f : errs =          63'b000000000000000000000000000000000000000000000000000000010010000; // D (0x0000000000000090) 
    12'ha03 : errs =          63'b000000000000000000000000000000000000000000000000000000010100000; // D (0x00000000000000a0) 
    12'hc02 : errs =          63'b000000000000000000000000000000000000000000000000000000011000000; // D (0x00000000000000c0) 
    12'h4eb : errs =          63'b000000000000000000000000000000000000000000000000000000010000000; // S (0x0000000000000080) 
//    12'hd3d : errs =          63'b000000000000000000000000000000000000000000000000000000110000000; // D (0x0000000000000180) 
//    12'h27e : errs =          63'b000000000000000000000000000000000000000000000000000001010000000; // D (0x0000000000000280) 
//    12'h9c1 : errs =          63'b000000000000000000000000000000000000000000000000000010010000000; // D (0x0000000000000480) 
//    12'hb86 : errs =          63'b000000000000000000000000000000000000000000000000000100010000000; // D (0x0000000000000880) 
//    12'hf08 : errs =          63'b000000000000000000000000000000000000000000000000001000010000000; // D (0x0000000000001080) 
//    12'h614 : errs =          63'b000000000000000000000000000000000000000000000000010000010000000; // D (0x0000000000002080) 
//    12'h115 : errs =          63'b000000000000000000000000000000000000000000000000100000010000000; // D (0x0000000000004080) 
//    12'hf17 : errs =          63'b000000000000000000000000000000000000000000000001000000010000000; // D (0x0000000000008080) 
//    12'h62a : errs =          63'b000000000000000000000000000000000000000000000010000000010000000; // D (0x0000000000010080) 
//    12'h169 : errs =          63'b000000000000000000000000000000000000000000000100000000010000000; // D (0x0000000000020080) 
//    12'hfef : errs =          63'b000000000000000000000000000000000000000000001000000000010000000; // D (0x0000000000040080) 
//    12'h7da : errs =          63'b000000000000000000000000000000000000000000010000000000010000000; // D (0x0000000000080080) 
//    12'h289 : errs =          63'b000000000000000000000000000000000000000000100000000000010000000; // D (0x0000000000100080) 
//    12'h82f : errs =          63'b000000000000000000000000000000000000000001000000000000010000000; // D (0x0000000000200080) 
//    12'h85a : errs =          63'b000000000000000000000000000000000000000010000000000000010000000; // D (0x0000000000400080) 
//    12'h8b0 : errs =          63'b000000000000000000000000000000000000000100000000000000010000000; // D (0x0000000000800080) 
//    12'h964 : errs =          63'b000000000000000000000000000000000000001000000000000000010000000; // D (0x0000000001000080) 
//    12'hacc : errs =          63'b000000000000000000000000000000000000010000000000000000010000000; // D (0x0000000002000080) 
//    12'hd9c : errs =          63'b000000000000000000000000000000000000100000000000000000010000000; // D (0x0000000004000080) 
//    12'h33c : errs =          63'b000000000000000000000000000000000001000000000000000000010000000; // D (0x0000000008000080) 
//    12'hb45 : errs =          63'b000000000000000000000000000000000010000000000000000000010000000; // D (0x0000000010000080) 
//    12'he8e : errs =          63'b000000000000000000000000000000000100000000000000000000010000000; // D (0x0000000020000080) 
//    12'h518 : errs =          63'b000000000000000000000000000000001000000000000000000000010000000; // D (0x0000000040000080) 
//    12'h70d : errs =          63'b000000000000000000000000000000010000000000000000000000010000000; // D (0x0000000080000080) 
//    12'h327 : errs =          63'b000000000000000000000000000000100000000000000000000000010000000; // D (0x0000000100000080) 
//    12'hb73 : errs =          63'b000000000000000000000000000001000000000000000000000000010000000; // D (0x0000000200000080) 
//    12'hee2 : errs =          63'b000000000000000000000000000010000000000000000000000000010000000; // D (0x0000000400000080) 
//    12'h5c0 : errs =          63'b000000000000000000000000000100000000000000000000000000010000000; // D (0x0000000800000080) 
//    12'h6bd : errs =          63'b000000000000000000000000001000000000000000000000000000010000000; // D (0x0000001000000080) 
//    12'h047 : errs =          63'b000000000000000000000000010000000000000000000000000000010000000; // D (0x0000002000000080) 
//    12'hdb3 : errs =          63'b000000000000000000000000100000000000000000000000000000010000000; // D (0x0000004000000080) 
//    12'h362 : errs =          63'b000000000000000000000001000000000000000000000000000000010000000; // D (0x0000008000000080) 
//    12'hbf9 : errs =          63'b000000000000000000000010000000000000000000000000000000010000000; // D (0x0000010000000080) 
//    12'hff6 : errs =          63'b000000000000000000000100000000000000000000000000000000010000000; // D (0x0000020000000080) 
//    12'h7e8 : errs =          63'b000000000000000000001000000000000000000000000000000000010000000; // D (0x0000040000000080) 
//    12'h2ed : errs =          63'b000000000000000000010000000000000000000000000000000000010000000; // D (0x0000080000000080) 
//    12'h8e7 : errs =          63'b000000000000000000100000000000000000000000000000000000010000000; // D (0x0000100000000080) 
//    12'h9ca : errs =          63'b000000000000000001000000000000000000000000000000000000010000000; // D (0x0000200000000080) 
//    12'hb90 : errs =          63'b000000000000000010000000000000000000000000000000000000010000000; // D (0x0000400000000080) 
//    12'hf24 : errs =          63'b000000000000000100000000000000000000000000000000000000010000000; // D (0x0000800000000080) 
//    12'h64c : errs =          63'b000000000000001000000000000000000000000000000000000000010000000; // D (0x0001000000000080) 
//    12'h1a5 : errs =          63'b000000000000010000000000000000000000000000000000000000010000000; // D (0x0002000000000080) 
//    12'he77 : errs =          63'b000000000000100000000000000000000000000000000000000000010000000; // D (0x0004000000000080) 
//    12'h4ea : errs =          63'b000000000001000000000000000000000000000000000000000000010000000; // D (0x0008000000000080) 
//    12'h4e9 : errs =          63'b000000000010000000000000000000000000000000000000000000010000000; // D (0x0010000000000080) 
//    12'h4ef : errs =          63'b000000000100000000000000000000000000000000000000000000010000000; // D (0x0020000000000080) 
//    12'h4e3 : errs =          63'b000000001000000000000000000000000000000000000000000000010000000; // D (0x0040000000000080) 
//    12'h4fb : errs =          63'b000000010000000000000000000000000000000000000000000000010000000; // D (0x0080000000000080) 
//    12'h4cb : errs =          63'b000000100000000000000000000000000000000000000000000000010000000; // D (0x0100000000000080) 
//    12'h4ab : errs =          63'b000001000000000000000000000000000000000000000000000000010000000; // D (0x0200000000000080) 
//    12'h46b : errs =          63'b000010000000000000000000000000000000000000000000000000010000000; // D (0x0400000000000080) 
//    12'h5eb : errs =          63'b000100000000000000000000000000000000000000000000000000010000000; // D (0x0800000000000080) 
//    12'h6eb : errs =          63'b001000000000000000000000000000000000000000000000000000010000000; // D (0x1000000000000080) 
//    12'h0eb : errs =          63'b010000000000000000000000000000000000000000000000000000010000000; // D (0x2000000000000080) 
//    12'hceb : errs =          63'b100000000000000000000000000000000000000000000000000000010000000; // D (0x4000000000000080) 
    12'hcef : errs =          63'b000000000000000000000000000000000000000000000000000000100000001; // D (0x0000000000000101) 
    12'h3a4 : errs =          63'b000000000000000000000000000000000000000000000000000000100000010; // D (0x0000000000000102) 
    12'h80b : errs =          63'b000000000000000000000000000000000000000000000000000000100000100; // D (0x0000000000000104) 
    12'ha6c : errs =          63'b000000000000000000000000000000000000000000000000000000100001000; // D (0x0000000000000108) 
    12'hea2 : errs =          63'b000000000000000000000000000000000000000000000000000000100010000; // D (0x0000000000000110) 
    12'h73e : errs =          63'b000000000000000000000000000000000000000000000000000000100100000; // D (0x0000000000000120) 
    12'h13f : errs =          63'b000000000000000000000000000000000000000000000000000000101000000; // D (0x0000000000000140) 
    12'hd3d : errs =          63'b000000000000000000000000000000000000000000000000000000110000000; // D (0x0000000000000180) 
    12'h9d6 : errs =          63'b000000000000000000000000000000000000000000000000000000100000000; // S (0x0000000000000100) 
//    12'hf43 : errs =          63'b000000000000000000000000000000000000000000000000000001100000000; // D (0x0000000000000300) 
//    12'h4fc : errs =          63'b000000000000000000000000000000000000000000000000000010100000000; // D (0x0000000000000500) 
//    12'h6bb : errs =          63'b000000000000000000000000000000000000000000000000000100100000000; // D (0x0000000000000900) 
//    12'h235 : errs =          63'b000000000000000000000000000000000000000000000000001000100000000; // D (0x0000000000001100) 
//    12'hb29 : errs =          63'b000000000000000000000000000000000000000000000000010000100000000; // D (0x0000000000002100) 
//    12'hc28 : errs =          63'b000000000000000000000000000000000000000000000000100000100000000; // D (0x0000000000004100) 
//    12'h22a : errs =          63'b000000000000000000000000000000000000000000000001000000100000000; // D (0x0000000000008100) 
//    12'hb17 : errs =          63'b000000000000000000000000000000000000000000000010000000100000000; // D (0x0000000000010100) 
//    12'hc54 : errs =          63'b000000000000000000000000000000000000000000000100000000100000000; // D (0x0000000000020100) 
//    12'h2d2 : errs =          63'b000000000000000000000000000000000000000000001000000000100000000; // D (0x0000000000040100) 
//    12'hae7 : errs =          63'b000000000000000000000000000000000000000000010000000000100000000; // D (0x0000000000080100) 
//    12'hfb4 : errs =          63'b000000000000000000000000000000000000000000100000000000100000000; // D (0x0000000000100100) 
//    12'h512 : errs =          63'b000000000000000000000000000000000000000001000000000000100000000; // D (0x0000000000200100) 
//    12'h567 : errs =          63'b000000000000000000000000000000000000000010000000000000100000000; // D (0x0000000000400100) 
//    12'h58d : errs =          63'b000000000000000000000000000000000000000100000000000000100000000; // D (0x0000000000800100) 
//    12'h459 : errs =          63'b000000000000000000000000000000000000001000000000000000100000000; // D (0x0000000001000100) 
//    12'h7f1 : errs =          63'b000000000000000000000000000000000000010000000000000000100000000; // D (0x0000000002000100) 
//    12'h0a1 : errs =          63'b000000000000000000000000000000000000100000000000000000100000000; // D (0x0000000004000100) 
//    12'he01 : errs =          63'b000000000000000000000000000000000001000000000000000000100000000; // D (0x0000000008000100) 
//    12'h678 : errs =          63'b000000000000000000000000000000000010000000000000000000100000000; // D (0x0000000010000100) 
//    12'h3b3 : errs =          63'b000000000000000000000000000000000100000000000000000000100000000; // D (0x0000000020000100) 
//    12'h825 : errs =          63'b000000000000000000000000000000001000000000000000000000100000000; // D (0x0000000040000100) 
//    12'ha30 : errs =          63'b000000000000000000000000000000010000000000000000000000100000000; // D (0x0000000080000100) 
//    12'he1a : errs =          63'b000000000000000000000000000000100000000000000000000000100000000; // D (0x0000000100000100) 
//    12'h64e : errs =          63'b000000000000000000000000000001000000000000000000000000100000000; // D (0x0000000200000100) 
//    12'h3df : errs =          63'b000000000000000000000000000010000000000000000000000000100000000; // D (0x0000000400000100) 
//    12'h8fd : errs =          63'b000000000000000000000000000100000000000000000000000000100000000; // D (0x0000000800000100) 
//    12'hb80 : errs =          63'b000000000000000000000000001000000000000000000000000000100000000; // D (0x0000001000000100) 
//    12'hd7a : errs =          63'b000000000000000000000000010000000000000000000000000000100000000; // D (0x0000002000000100) 
//    12'h08e : errs =          63'b000000000000000000000000100000000000000000000000000000100000000; // D (0x0000004000000100) 
//    12'he5f : errs =          63'b000000000000000000000001000000000000000000000000000000100000000; // D (0x0000008000000100) 
//    12'h6c4 : errs =          63'b000000000000000000000010000000000000000000000000000000100000000; // D (0x0000010000000100) 
//    12'h2cb : errs =          63'b000000000000000000000100000000000000000000000000000000100000000; // D (0x0000020000000100) 
//    12'had5 : errs =          63'b000000000000000000001000000000000000000000000000000000100000000; // D (0x0000040000000100) 
//    12'hfd0 : errs =          63'b000000000000000000010000000000000000000000000000000000100000000; // D (0x0000080000000100) 
//    12'h5da : errs =          63'b000000000000000000100000000000000000000000000000000000100000000; // D (0x0000100000000100) 
//    12'h4f7 : errs =          63'b000000000000000001000000000000000000000000000000000000100000000; // D (0x0000200000000100) 
//    12'h6ad : errs =          63'b000000000000000010000000000000000000000000000000000000100000000; // D (0x0000400000000100) 
//    12'h219 : errs =          63'b000000000000000100000000000000000000000000000000000000100000000; // D (0x0000800000000100) 
//    12'hb71 : errs =          63'b000000000000001000000000000000000000000000000000000000100000000; // D (0x0001000000000100) 
//    12'hc98 : errs =          63'b000000000000010000000000000000000000000000000000000000100000000; // D (0x0002000000000100) 
//    12'h34a : errs =          63'b000000000000100000000000000000000000000000000000000000100000000; // D (0x0004000000000100) 
//    12'h9d7 : errs =          63'b000000000001000000000000000000000000000000000000000000100000000; // D (0x0008000000000100) 
//    12'h9d4 : errs =          63'b000000000010000000000000000000000000000000000000000000100000000; // D (0x0010000000000100) 
//    12'h9d2 : errs =          63'b000000000100000000000000000000000000000000000000000000100000000; // D (0x0020000000000100) 
//    12'h9de : errs =          63'b000000001000000000000000000000000000000000000000000000100000000; // D (0x0040000000000100) 
//    12'h9c6 : errs =          63'b000000010000000000000000000000000000000000000000000000100000000; // D (0x0080000000000100) 
//    12'h9f6 : errs =          63'b000000100000000000000000000000000000000000000000000000100000000; // D (0x0100000000000100) 
//    12'h996 : errs =          63'b000001000000000000000000000000000000000000000000000000100000000; // D (0x0200000000000100) 
//    12'h956 : errs =          63'b000010000000000000000000000000000000000000000000000000100000000; // D (0x0400000000000100) 
//    12'h8d6 : errs =          63'b000100000000000000000000000000000000000000000000000000100000000; // D (0x0800000000000100) 
//    12'hbd6 : errs =          63'b001000000000000000000000000000000000000000000000000000100000000; // D (0x1000000000000100) 
//    12'hdd6 : errs =          63'b010000000000000000000000000000000000000000000000000000100000000; // D (0x2000000000000100) 
//    12'h1d6 : errs =          63'b100000000000000000000000000000000000000000000000000000100000000; // D (0x4000000000000100) 
    12'h3ac : errs =          63'b000000000000000000000000000000000000000000000000000001000000001; // D (0x0000000000000201) 
    12'hce7 : errs =          63'b000000000000000000000000000000000000000000000000000001000000010; // D (0x0000000000000202) 
    12'h748 : errs =          63'b000000000000000000000000000000000000000000000000000001000000100; // D (0x0000000000000204) 
    12'h52f : errs =          63'b000000000000000000000000000000000000000000000000000001000001000; // D (0x0000000000000208) 
    12'h1e1 : errs =          63'b000000000000000000000000000000000000000000000000000001000010000; // D (0x0000000000000210) 
    12'h87d : errs =          63'b000000000000000000000000000000000000000000000000000001000100000; // D (0x0000000000000220) 
    12'he7c : errs =          63'b000000000000000000000000000000000000000000000000000001001000000; // D (0x0000000000000240) 
    12'h27e : errs =          63'b000000000000000000000000000000000000000000000000000001010000000; // D (0x0000000000000280) 
    12'hf43 : errs =          63'b000000000000000000000000000000000000000000000000000001100000000; // D (0x0000000000000300) 
    12'h695 : errs =          63'b000000000000000000000000000000000000000000000000000001000000000; // S (0x0000000000000200) 
//    12'hbbf : errs =          63'b000000000000000000000000000000000000000000000000000011000000000; // D (0x0000000000000600) 
//    12'h9f8 : errs =          63'b000000000000000000000000000000000000000000000000000101000000000; // D (0x0000000000000a00) 
//    12'hd76 : errs =          63'b000000000000000000000000000000000000000000000000001001000000000; // D (0x0000000000001200) 
//    12'h46a : errs =          63'b000000000000000000000000000000000000000000000000010001000000000; // D (0x0000000000002200) 
//    12'h36b : errs =          63'b000000000000000000000000000000000000000000000000100001000000000; // D (0x0000000000004200) 
//    12'hd69 : errs =          63'b000000000000000000000000000000000000000000000001000001000000000; // D (0x0000000000008200) 
//    12'h454 : errs =          63'b000000000000000000000000000000000000000000000010000001000000000; // D (0x0000000000010200) 
//    12'h317 : errs =          63'b000000000000000000000000000000000000000000000100000001000000000; // D (0x0000000000020200) 
//    12'hd91 : errs =          63'b000000000000000000000000000000000000000000001000000001000000000; // D (0x0000000000040200) 
//    12'h5a4 : errs =          63'b000000000000000000000000000000000000000000010000000001000000000; // D (0x0000000000080200) 
//    12'h0f7 : errs =          63'b000000000000000000000000000000000000000000100000000001000000000; // D (0x0000000000100200) 
//    12'ha51 : errs =          63'b000000000000000000000000000000000000000001000000000001000000000; // D (0x0000000000200200) 
//    12'ha24 : errs =          63'b000000000000000000000000000000000000000010000000000001000000000; // D (0x0000000000400200) 
//    12'hace : errs =          63'b000000000000000000000000000000000000000100000000000001000000000; // D (0x0000000000800200) 
//    12'hb1a : errs =          63'b000000000000000000000000000000000000001000000000000001000000000; // D (0x0000000001000200) 
//    12'h8b2 : errs =          63'b000000000000000000000000000000000000010000000000000001000000000; // D (0x0000000002000200) 
//    12'hfe2 : errs =          63'b000000000000000000000000000000000000100000000000000001000000000; // D (0x0000000004000200) 
//    12'h142 : errs =          63'b000000000000000000000000000000000001000000000000000001000000000; // D (0x0000000008000200) 
//    12'h93b : errs =          63'b000000000000000000000000000000000010000000000000000001000000000; // D (0x0000000010000200) 
//    12'hcf0 : errs =          63'b000000000000000000000000000000000100000000000000000001000000000; // D (0x0000000020000200) 
//    12'h766 : errs =          63'b000000000000000000000000000000001000000000000000000001000000000; // D (0x0000000040000200) 
//    12'h573 : errs =          63'b000000000000000000000000000000010000000000000000000001000000000; // D (0x0000000080000200) 
//    12'h159 : errs =          63'b000000000000000000000000000000100000000000000000000001000000000; // D (0x0000000100000200) 
//    12'h90d : errs =          63'b000000000000000000000000000001000000000000000000000001000000000; // D (0x0000000200000200) 
//    12'hc9c : errs =          63'b000000000000000000000000000010000000000000000000000001000000000; // D (0x0000000400000200) 
//    12'h7be : errs =          63'b000000000000000000000000000100000000000000000000000001000000000; // D (0x0000000800000200) 
//    12'h4c3 : errs =          63'b000000000000000000000000001000000000000000000000000001000000000; // D (0x0000001000000200) 
//    12'h239 : errs =          63'b000000000000000000000000010000000000000000000000000001000000000; // D (0x0000002000000200) 
//    12'hfcd : errs =          63'b000000000000000000000000100000000000000000000000000001000000000; // D (0x0000004000000200) 
//    12'h11c : errs =          63'b000000000000000000000001000000000000000000000000000001000000000; // D (0x0000008000000200) 
//    12'h987 : errs =          63'b000000000000000000000010000000000000000000000000000001000000000; // D (0x0000010000000200) 
//    12'hd88 : errs =          63'b000000000000000000000100000000000000000000000000000001000000000; // D (0x0000020000000200) 
//    12'h596 : errs =          63'b000000000000000000001000000000000000000000000000000001000000000; // D (0x0000040000000200) 
//    12'h093 : errs =          63'b000000000000000000010000000000000000000000000000000001000000000; // D (0x0000080000000200) 
//    12'ha99 : errs =          63'b000000000000000000100000000000000000000000000000000001000000000; // D (0x0000100000000200) 
//    12'hbb4 : errs =          63'b000000000000000001000000000000000000000000000000000001000000000; // D (0x0000200000000200) 
//    12'h9ee : errs =          63'b000000000000000010000000000000000000000000000000000001000000000; // D (0x0000400000000200) 
//    12'hd5a : errs =          63'b000000000000000100000000000000000000000000000000000001000000000; // D (0x0000800000000200) 
//    12'h432 : errs =          63'b000000000000001000000000000000000000000000000000000001000000000; // D (0x0001000000000200) 
//    12'h3db : errs =          63'b000000000000010000000000000000000000000000000000000001000000000; // D (0x0002000000000200) 
//    12'hc09 : errs =          63'b000000000000100000000000000000000000000000000000000001000000000; // D (0x0004000000000200) 
//    12'h694 : errs =          63'b000000000001000000000000000000000000000000000000000001000000000; // D (0x0008000000000200) 
//    12'h697 : errs =          63'b000000000010000000000000000000000000000000000000000001000000000; // D (0x0010000000000200) 
//    12'h691 : errs =          63'b000000000100000000000000000000000000000000000000000001000000000; // D (0x0020000000000200) 
//    12'h69d : errs =          63'b000000001000000000000000000000000000000000000000000001000000000; // D (0x0040000000000200) 
//    12'h685 : errs =          63'b000000010000000000000000000000000000000000000000000001000000000; // D (0x0080000000000200) 
//    12'h6b5 : errs =          63'b000000100000000000000000000000000000000000000000000001000000000; // D (0x0100000000000200) 
//    12'h6d5 : errs =          63'b000001000000000000000000000000000000000000000000000001000000000; // D (0x0200000000000200) 
//    12'h615 : errs =          63'b000010000000000000000000000000000000000000000000000001000000000; // D (0x0400000000000200) 
//    12'h795 : errs =          63'b000100000000000000000000000000000000000000000000000001000000000; // D (0x0800000000000200) 
//    12'h495 : errs =          63'b001000000000000000000000000000000000000000000000000001000000000; // D (0x1000000000000200) 
//    12'h295 : errs =          63'b010000000000000000000000000000000000000000000000000001000000000; // D (0x2000000000000200) 
//    12'he95 : errs =          63'b100000000000000000000000000000000000000000000000000001000000000; // D (0x4000000000000200) 
    12'h813 : errs =          63'b000000000000000000000000000000000000000000000000000010000000001; // D (0x0000000000000401) 
    12'h758 : errs =          63'b000000000000000000000000000000000000000000000000000010000000010; // D (0x0000000000000402) 
    12'hcf7 : errs =          63'b000000000000000000000000000000000000000000000000000010000000100; // D (0x0000000000000404) 
    12'he90 : errs =          63'b000000000000000000000000000000000000000000000000000010000001000; // D (0x0000000000000408) 
    12'ha5e : errs =          63'b000000000000000000000000000000000000000000000000000010000010000; // D (0x0000000000000410) 
    12'h3c2 : errs =          63'b000000000000000000000000000000000000000000000000000010000100000; // D (0x0000000000000420) 
    12'h5c3 : errs =          63'b000000000000000000000000000000000000000000000000000010001000000; // D (0x0000000000000440) 
    12'h9c1 : errs =          63'b000000000000000000000000000000000000000000000000000010010000000; // D (0x0000000000000480) 
    12'h4fc : errs =          63'b000000000000000000000000000000000000000000000000000010100000000; // D (0x0000000000000500) 
    12'hbbf : errs =          63'b000000000000000000000000000000000000000000000000000011000000000; // D (0x0000000000000600) 
    12'hd2a : errs =          63'b000000000000000000000000000000000000000000000000000010000000000; // S (0x0000000000000400) 
//    12'h247 : errs =          63'b000000000000000000000000000000000000000000000000000110000000000; // D (0x0000000000000c00) 
//    12'h6c9 : errs =          63'b000000000000000000000000000000000000000000000000001010000000000; // D (0x0000000000001400) 
//    12'hfd5 : errs =          63'b000000000000000000000000000000000000000000000000010010000000000; // D (0x0000000000002400) 
//    12'h8d4 : errs =          63'b000000000000000000000000000000000000000000000000100010000000000; // D (0x0000000000004400) 
//    12'h6d6 : errs =          63'b000000000000000000000000000000000000000000000001000010000000000; // D (0x0000000000008400) 
//    12'hfeb : errs =          63'b000000000000000000000000000000000000000000000010000010000000000; // D (0x0000000000010400) 
//    12'h8a8 : errs =          63'b000000000000000000000000000000000000000000000100000010000000000; // D (0x0000000000020400) 
//    12'h62e : errs =          63'b000000000000000000000000000000000000000000001000000010000000000; // D (0x0000000000040400) 
//    12'he1b : errs =          63'b000000000000000000000000000000000000000000010000000010000000000; // D (0x0000000000080400) 
//    12'hb48 : errs =          63'b000000000000000000000000000000000000000000100000000010000000000; // D (0x0000000000100400) 
//    12'h1ee : errs =          63'b000000000000000000000000000000000000000001000000000010000000000; // D (0x0000000000200400) 
//    12'h19b : errs =          63'b000000000000000000000000000000000000000010000000000010000000000; // D (0x0000000000400400) 
//    12'h171 : errs =          63'b000000000000000000000000000000000000000100000000000010000000000; // D (0x0000000000800400) 
//    12'h0a5 : errs =          63'b000000000000000000000000000000000000001000000000000010000000000; // D (0x0000000001000400) 
//    12'h30d : errs =          63'b000000000000000000000000000000000000010000000000000010000000000; // D (0x0000000002000400) 
//    12'h45d : errs =          63'b000000000000000000000000000000000000100000000000000010000000000; // D (0x0000000004000400) 
//    12'hafd : errs =          63'b000000000000000000000000000000000001000000000000000010000000000; // D (0x0000000008000400) 
//    12'h284 : errs =          63'b000000000000000000000000000000000010000000000000000010000000000; // D (0x0000000010000400) 
//    12'h74f : errs =          63'b000000000000000000000000000000000100000000000000000010000000000; // D (0x0000000020000400) 
//    12'hcd9 : errs =          63'b000000000000000000000000000000001000000000000000000010000000000; // D (0x0000000040000400) 
//    12'hecc : errs =          63'b000000000000000000000000000000010000000000000000000010000000000; // D (0x0000000080000400) 
//    12'hae6 : errs =          63'b000000000000000000000000000000100000000000000000000010000000000; // D (0x0000000100000400) 
//    12'h2b2 : errs =          63'b000000000000000000000000000001000000000000000000000010000000000; // D (0x0000000200000400) 
//    12'h723 : errs =          63'b000000000000000000000000000010000000000000000000000010000000000; // D (0x0000000400000400) 
//    12'hc01 : errs =          63'b000000000000000000000000000100000000000000000000000010000000000; // D (0x0000000800000400) 
//    12'hf7c : errs =          63'b000000000000000000000000001000000000000000000000000010000000000; // D (0x0000001000000400) 
//    12'h986 : errs =          63'b000000000000000000000000010000000000000000000000000010000000000; // D (0x0000002000000400) 
//    12'h472 : errs =          63'b000000000000000000000000100000000000000000000000000010000000000; // D (0x0000004000000400) 
//    12'haa3 : errs =          63'b000000000000000000000001000000000000000000000000000010000000000; // D (0x0000008000000400) 
//    12'h238 : errs =          63'b000000000000000000000010000000000000000000000000000010000000000; // D (0x0000010000000400) 
//    12'h637 : errs =          63'b000000000000000000000100000000000000000000000000000010000000000; // D (0x0000020000000400) 
//    12'he29 : errs =          63'b000000000000000000001000000000000000000000000000000010000000000; // D (0x0000040000000400) 
//    12'hb2c : errs =          63'b000000000000000000010000000000000000000000000000000010000000000; // D (0x0000080000000400) 
//    12'h126 : errs =          63'b000000000000000000100000000000000000000000000000000010000000000; // D (0x0000100000000400) 
//    12'h00b : errs =          63'b000000000000000001000000000000000000000000000000000010000000000; // D (0x0000200000000400) 
//    12'h251 : errs =          63'b000000000000000010000000000000000000000000000000000010000000000; // D (0x0000400000000400) 
//    12'h6e5 : errs =          63'b000000000000000100000000000000000000000000000000000010000000000; // D (0x0000800000000400) 
//    12'hf8d : errs =          63'b000000000000001000000000000000000000000000000000000010000000000; // D (0x0001000000000400) 
//    12'h864 : errs =          63'b000000000000010000000000000000000000000000000000000010000000000; // D (0x0002000000000400) 
//    12'h7b6 : errs =          63'b000000000000100000000000000000000000000000000000000010000000000; // D (0x0004000000000400) 
//    12'hd2b : errs =          63'b000000000001000000000000000000000000000000000000000010000000000; // D (0x0008000000000400) 
//    12'hd28 : errs =          63'b000000000010000000000000000000000000000000000000000010000000000; // D (0x0010000000000400) 
//    12'hd2e : errs =          63'b000000000100000000000000000000000000000000000000000010000000000; // D (0x0020000000000400) 
//    12'hd22 : errs =          63'b000000001000000000000000000000000000000000000000000010000000000; // D (0x0040000000000400) 
//    12'hd3a : errs =          63'b000000010000000000000000000000000000000000000000000010000000000; // D (0x0080000000000400) 
//    12'hd0a : errs =          63'b000000100000000000000000000000000000000000000000000010000000000; // D (0x0100000000000400) 
//    12'hd6a : errs =          63'b000001000000000000000000000000000000000000000000000010000000000; // D (0x0200000000000400) 
//    12'hdaa : errs =          63'b000010000000000000000000000000000000000000000000000010000000000; // D (0x0400000000000400) 
//    12'hc2a : errs =          63'b000100000000000000000000000000000000000000000000000010000000000; // D (0x0800000000000400) 
//    12'hf2a : errs =          63'b001000000000000000000000000000000000000000000000000010000000000; // D (0x1000000000000400) 
//    12'h92a : errs =          63'b010000000000000000000000000000000000000000000000000010000000000; // D (0x2000000000000400) 
//    12'h52a : errs =          63'b100000000000000000000000000000000000000000000000000010000000000; // D (0x4000000000000400) 
    12'ha54 : errs =          63'b000000000000000000000000000000000000000000000000000100000000001; // D (0x0000000000000801) 
    12'h51f : errs =          63'b000000000000000000000000000000000000000000000000000100000000010; // D (0x0000000000000802) 
    12'heb0 : errs =          63'b000000000000000000000000000000000000000000000000000100000000100; // D (0x0000000000000804) 
    12'hcd7 : errs =          63'b000000000000000000000000000000000000000000000000000100000001000; // D (0x0000000000000808) 
    12'h819 : errs =          63'b000000000000000000000000000000000000000000000000000100000010000; // D (0x0000000000000810) 
    12'h185 : errs =          63'b000000000000000000000000000000000000000000000000000100000100000; // D (0x0000000000000820) 
    12'h784 : errs =          63'b000000000000000000000000000000000000000000000000000100001000000; // D (0x0000000000000840) 
    12'hb86 : errs =          63'b000000000000000000000000000000000000000000000000000100010000000; // D (0x0000000000000880) 
    12'h6bb : errs =          63'b000000000000000000000000000000000000000000000000000100100000000; // D (0x0000000000000900) 
    12'h9f8 : errs =          63'b000000000000000000000000000000000000000000000000000101000000000; // D (0x0000000000000a00) 
    12'h247 : errs =          63'b000000000000000000000000000000000000000000000000000110000000000; // D (0x0000000000000c00) 
    12'hf6d : errs =          63'b000000000000000000000000000000000000000000000000000100000000000; // S (0x0000000000000800) 
//    12'h48e : errs =          63'b000000000000000000000000000000000000000000000000001100000000000; // D (0x0000000000001800) 
//    12'hd92 : errs =          63'b000000000000000000000000000000000000000000000000010100000000000; // D (0x0000000000002800) 
//    12'ha93 : errs =          63'b000000000000000000000000000000000000000000000000100100000000000; // D (0x0000000000004800) 
//    12'h491 : errs =          63'b000000000000000000000000000000000000000000000001000100000000000; // D (0x0000000000008800) 
//    12'hdac : errs =          63'b000000000000000000000000000000000000000000000010000100000000000; // D (0x0000000000010800) 
//    12'haef : errs =          63'b000000000000000000000000000000000000000000000100000100000000000; // D (0x0000000000020800) 
//    12'h469 : errs =          63'b000000000000000000000000000000000000000000001000000100000000000; // D (0x0000000000040800) 
//    12'hc5c : errs =          63'b000000000000000000000000000000000000000000010000000100000000000; // D (0x0000000000080800) 
//    12'h90f : errs =          63'b000000000000000000000000000000000000000000100000000100000000000; // D (0x0000000000100800) 
//    12'h3a9 : errs =          63'b000000000000000000000000000000000000000001000000000100000000000; // D (0x0000000000200800) 
//    12'h3dc : errs =          63'b000000000000000000000000000000000000000010000000000100000000000; // D (0x0000000000400800) 
//    12'h336 : errs =          63'b000000000000000000000000000000000000000100000000000100000000000; // D (0x0000000000800800) 
//    12'h2e2 : errs =          63'b000000000000000000000000000000000000001000000000000100000000000; // D (0x0000000001000800) 
//    12'h14a : errs =          63'b000000000000000000000000000000000000010000000000000100000000000; // D (0x0000000002000800) 
//    12'h61a : errs =          63'b000000000000000000000000000000000000100000000000000100000000000; // D (0x0000000004000800) 
//    12'h8ba : errs =          63'b000000000000000000000000000000000001000000000000000100000000000; // D (0x0000000008000800) 
//    12'h0c3 : errs =          63'b000000000000000000000000000000000010000000000000000100000000000; // D (0x0000000010000800) 
//    12'h508 : errs =          63'b000000000000000000000000000000000100000000000000000100000000000; // D (0x0000000020000800) 
//    12'he9e : errs =          63'b000000000000000000000000000000001000000000000000000100000000000; // D (0x0000000040000800) 
//    12'hc8b : errs =          63'b000000000000000000000000000000010000000000000000000100000000000; // D (0x0000000080000800) 
//    12'h8a1 : errs =          63'b000000000000000000000000000000100000000000000000000100000000000; // D (0x0000000100000800) 
//    12'h0f5 : errs =          63'b000000000000000000000000000001000000000000000000000100000000000; // D (0x0000000200000800) 
//    12'h564 : errs =          63'b000000000000000000000000000010000000000000000000000100000000000; // D (0x0000000400000800) 
//    12'he46 : errs =          63'b000000000000000000000000000100000000000000000000000100000000000; // D (0x0000000800000800) 
//    12'hd3b : errs =          63'b000000000000000000000000001000000000000000000000000100000000000; // D (0x0000001000000800) 
//    12'hbc1 : errs =          63'b000000000000000000000000010000000000000000000000000100000000000; // D (0x0000002000000800) 
//    12'h635 : errs =          63'b000000000000000000000000100000000000000000000000000100000000000; // D (0x0000004000000800) 
//    12'h8e4 : errs =          63'b000000000000000000000001000000000000000000000000000100000000000; // D (0x0000008000000800) 
//    12'h07f : errs =          63'b000000000000000000000010000000000000000000000000000100000000000; // D (0x0000010000000800) 
//    12'h470 : errs =          63'b000000000000000000000100000000000000000000000000000100000000000; // D (0x0000020000000800) 
//    12'hc6e : errs =          63'b000000000000000000001000000000000000000000000000000100000000000; // D (0x0000040000000800) 
//    12'h96b : errs =          63'b000000000000000000010000000000000000000000000000000100000000000; // D (0x0000080000000800) 
//    12'h361 : errs =          63'b000000000000000000100000000000000000000000000000000100000000000; // D (0x0000100000000800) 
//    12'h24c : errs =          63'b000000000000000001000000000000000000000000000000000100000000000; // D (0x0000200000000800) 
//    12'h016 : errs =          63'b000000000000000010000000000000000000000000000000000100000000000; // D (0x0000400000000800) 
//    12'h4a2 : errs =          63'b000000000000000100000000000000000000000000000000000100000000000; // D (0x0000800000000800) 
//    12'hdca : errs =          63'b000000000000001000000000000000000000000000000000000100000000000; // D (0x0001000000000800) 
//    12'ha23 : errs =          63'b000000000000010000000000000000000000000000000000000100000000000; // D (0x0002000000000800) 
//    12'h5f1 : errs =          63'b000000000000100000000000000000000000000000000000000100000000000; // D (0x0004000000000800) 
//    12'hf6c : errs =          63'b000000000001000000000000000000000000000000000000000100000000000; // D (0x0008000000000800) 
//    12'hf6f : errs =          63'b000000000010000000000000000000000000000000000000000100000000000; // D (0x0010000000000800) 
//    12'hf69 : errs =          63'b000000000100000000000000000000000000000000000000000100000000000; // D (0x0020000000000800) 
//    12'hf65 : errs =          63'b000000001000000000000000000000000000000000000000000100000000000; // D (0x0040000000000800) 
//    12'hf7d : errs =          63'b000000010000000000000000000000000000000000000000000100000000000; // D (0x0080000000000800) 
//    12'hf4d : errs =          63'b000000100000000000000000000000000000000000000000000100000000000; // D (0x0100000000000800) 
//    12'hf2d : errs =          63'b000001000000000000000000000000000000000000000000000100000000000; // D (0x0200000000000800) 
//    12'hfed : errs =          63'b000010000000000000000000000000000000000000000000000100000000000; // D (0x0400000000000800) 
//    12'he6d : errs =          63'b000100000000000000000000000000000000000000000000000100000000000; // D (0x0800000000000800) 
//    12'hd6d : errs =          63'b001000000000000000000000000000000000000000000000000100000000000; // D (0x1000000000000800) 
//    12'hb6d : errs =          63'b010000000000000000000000000000000000000000000000000100000000000; // D (0x2000000000000800) 
//    12'h76d : errs =          63'b100000000000000000000000000000000000000000000000000100000000000; // D (0x4000000000000800) 
    12'heda : errs =          63'b000000000000000000000000000000000000000000000000001000000000001; // D (0x0000000000001001) 
    12'h191 : errs =          63'b000000000000000000000000000000000000000000000000001000000000010; // D (0x0000000000001002) 
    12'ha3e : errs =          63'b000000000000000000000000000000000000000000000000001000000000100; // D (0x0000000000001004) 
    12'h859 : errs =          63'b000000000000000000000000000000000000000000000000001000000001000; // D (0x0000000000001008) 
    12'hc97 : errs =          63'b000000000000000000000000000000000000000000000000001000000010000; // D (0x0000000000001010) 
    12'h50b : errs =          63'b000000000000000000000000000000000000000000000000001000000100000; // D (0x0000000000001020) 
    12'h30a : errs =          63'b000000000000000000000000000000000000000000000000001000001000000; // D (0x0000000000001040) 
    12'hf08 : errs =          63'b000000000000000000000000000000000000000000000000001000010000000; // D (0x0000000000001080) 
    12'h235 : errs =          63'b000000000000000000000000000000000000000000000000001000100000000; // D (0x0000000000001100) 
    12'hd76 : errs =          63'b000000000000000000000000000000000000000000000000001001000000000; // D (0x0000000000001200) 
    12'h6c9 : errs =          63'b000000000000000000000000000000000000000000000000001010000000000; // D (0x0000000000001400) 
    12'h48e : errs =          63'b000000000000000000000000000000000000000000000000001100000000000; // D (0x0000000000001800) 
    12'hbe3 : errs =          63'b000000000000000000000000000000000000000000000000001000000000000; // S (0x0000000000001000) 
//    12'h91c : errs =          63'b000000000000000000000000000000000000000000000000011000000000000; // D (0x0000000000003000) 
//    12'he1d : errs =          63'b000000000000000000000000000000000000000000000000101000000000000; // D (0x0000000000005000) 
//    12'h01f : errs =          63'b000000000000000000000000000000000000000000000001001000000000000; // D (0x0000000000009000) 
//    12'h922 : errs =          63'b000000000000000000000000000000000000000000000010001000000000000; // D (0x0000000000011000) 
//    12'he61 : errs =          63'b000000000000000000000000000000000000000000000100001000000000000; // D (0x0000000000021000) 
//    12'h0e7 : errs =          63'b000000000000000000000000000000000000000000001000001000000000000; // D (0x0000000000041000) 
//    12'h8d2 : errs =          63'b000000000000000000000000000000000000000000010000001000000000000; // D (0x0000000000081000) 
//    12'hd81 : errs =          63'b000000000000000000000000000000000000000000100000001000000000000; // D (0x0000000000101000) 
//    12'h727 : errs =          63'b000000000000000000000000000000000000000001000000001000000000000; // D (0x0000000000201000) 
//    12'h752 : errs =          63'b000000000000000000000000000000000000000010000000001000000000000; // D (0x0000000000401000) 
//    12'h7b8 : errs =          63'b000000000000000000000000000000000000000100000000001000000000000; // D (0x0000000000801000) 
//    12'h66c : errs =          63'b000000000000000000000000000000000000001000000000001000000000000; // D (0x0000000001001000) 
//    12'h5c4 : errs =          63'b000000000000000000000000000000000000010000000000001000000000000; // D (0x0000000002001000) 
//    12'h294 : errs =          63'b000000000000000000000000000000000000100000000000001000000000000; // D (0x0000000004001000) 
//    12'hc34 : errs =          63'b000000000000000000000000000000000001000000000000001000000000000; // D (0x0000000008001000) 
//    12'h44d : errs =          63'b000000000000000000000000000000000010000000000000001000000000000; // D (0x0000000010001000) 
//    12'h186 : errs =          63'b000000000000000000000000000000000100000000000000001000000000000; // D (0x0000000020001000) 
//    12'ha10 : errs =          63'b000000000000000000000000000000001000000000000000001000000000000; // D (0x0000000040001000) 
//    12'h805 : errs =          63'b000000000000000000000000000000010000000000000000001000000000000; // D (0x0000000080001000) 
//    12'hc2f : errs =          63'b000000000000000000000000000000100000000000000000001000000000000; // D (0x0000000100001000) 
//    12'h47b : errs =          63'b000000000000000000000000000001000000000000000000001000000000000; // D (0x0000000200001000) 
//    12'h1ea : errs =          63'b000000000000000000000000000010000000000000000000001000000000000; // D (0x0000000400001000) 
//    12'hac8 : errs =          63'b000000000000000000000000000100000000000000000000001000000000000; // D (0x0000000800001000) 
//    12'h9b5 : errs =          63'b000000000000000000000000001000000000000000000000001000000000000; // D (0x0000001000001000) 
//    12'hf4f : errs =          63'b000000000000000000000000010000000000000000000000001000000000000; // D (0x0000002000001000) 
//    12'h2bb : errs =          63'b000000000000000000000000100000000000000000000000001000000000000; // D (0x0000004000001000) 
//    12'hc6a : errs =          63'b000000000000000000000001000000000000000000000000001000000000000; // D (0x0000008000001000) 
//    12'h4f1 : errs =          63'b000000000000000000000010000000000000000000000000001000000000000; // D (0x0000010000001000) 
//    12'h0fe : errs =          63'b000000000000000000000100000000000000000000000000001000000000000; // D (0x0000020000001000) 
//    12'h8e0 : errs =          63'b000000000000000000001000000000000000000000000000001000000000000; // D (0x0000040000001000) 
//    12'hde5 : errs =          63'b000000000000000000010000000000000000000000000000001000000000000; // D (0x0000080000001000) 
//    12'h7ef : errs =          63'b000000000000000000100000000000000000000000000000001000000000000; // D (0x0000100000001000) 
//    12'h6c2 : errs =          63'b000000000000000001000000000000000000000000000000001000000000000; // D (0x0000200000001000) 
//    12'h498 : errs =          63'b000000000000000010000000000000000000000000000000001000000000000; // D (0x0000400000001000) 
//    12'h02c : errs =          63'b000000000000000100000000000000000000000000000000001000000000000; // D (0x0000800000001000) 
//    12'h944 : errs =          63'b000000000000001000000000000000000000000000000000001000000000000; // D (0x0001000000001000) 
//    12'head : errs =          63'b000000000000010000000000000000000000000000000000001000000000000; // D (0x0002000000001000) 
//    12'h17f : errs =          63'b000000000000100000000000000000000000000000000000001000000000000; // D (0x0004000000001000) 
//    12'hbe2 : errs =          63'b000000000001000000000000000000000000000000000000001000000000000; // D (0x0008000000001000) 
//    12'hbe1 : errs =          63'b000000000010000000000000000000000000000000000000001000000000000; // D (0x0010000000001000) 
//    12'hbe7 : errs =          63'b000000000100000000000000000000000000000000000000001000000000000; // D (0x0020000000001000) 
//    12'hbeb : errs =          63'b000000001000000000000000000000000000000000000000001000000000000; // D (0x0040000000001000) 
//    12'hbf3 : errs =          63'b000000010000000000000000000000000000000000000000001000000000000; // D (0x0080000000001000) 
//    12'hbc3 : errs =          63'b000000100000000000000000000000000000000000000000001000000000000; // D (0x0100000000001000) 
//    12'hba3 : errs =          63'b000001000000000000000000000000000000000000000000001000000000000; // D (0x0200000000001000) 
//    12'hb63 : errs =          63'b000010000000000000000000000000000000000000000000001000000000000; // D (0x0400000000001000) 
//    12'hae3 : errs =          63'b000100000000000000000000000000000000000000000000001000000000000; // D (0x0800000000001000) 
//    12'h9e3 : errs =          63'b001000000000000000000000000000000000000000000000001000000000000; // D (0x1000000000001000) 
//    12'hfe3 : errs =          63'b010000000000000000000000000000000000000000000000001000000000000; // D (0x2000000000001000) 
//    12'h3e3 : errs =          63'b100000000000000000000000000000000000000000000000001000000000000; // D (0x4000000000001000) 
    12'h7c6 : errs =          63'b000000000000000000000000000000000000000000000000010000000000001; // D (0x0000000000002001) 
    12'h88d : errs =          63'b000000000000000000000000000000000000000000000000010000000000010; // D (0x0000000000002002) 
    12'h322 : errs =          63'b000000000000000000000000000000000000000000000000010000000000100; // D (0x0000000000002004) 
    12'h145 : errs =          63'b000000000000000000000000000000000000000000000000010000000001000; // D (0x0000000000002008) 
    12'h58b : errs =          63'b000000000000000000000000000000000000000000000000010000000010000; // D (0x0000000000002010) 
    12'hc17 : errs =          63'b000000000000000000000000000000000000000000000000010000000100000; // D (0x0000000000002020) 
    12'ha16 : errs =          63'b000000000000000000000000000000000000000000000000010000001000000; // D (0x0000000000002040) 
    12'h614 : errs =          63'b000000000000000000000000000000000000000000000000010000010000000; // D (0x0000000000002080) 
    12'hb29 : errs =          63'b000000000000000000000000000000000000000000000000010000100000000; // D (0x0000000000002100) 
    12'h46a : errs =          63'b000000000000000000000000000000000000000000000000010001000000000; // D (0x0000000000002200) 
    12'hfd5 : errs =          63'b000000000000000000000000000000000000000000000000010010000000000; // D (0x0000000000002400) 
    12'hd92 : errs =          63'b000000000000000000000000000000000000000000000000010100000000000; // D (0x0000000000002800) 
    12'h91c : errs =          63'b000000000000000000000000000000000000000000000000011000000000000; // D (0x0000000000003000) 
    12'h2ff : errs =          63'b000000000000000000000000000000000000000000000000010000000000000; // S (0x0000000000002000) 
//    12'h701 : errs =          63'b000000000000000000000000000000000000000000000000110000000000000; // D (0x0000000000006000) 
//    12'h903 : errs =          63'b000000000000000000000000000000000000000000000001010000000000000; // D (0x000000000000a000) 
//    12'h03e : errs =          63'b000000000000000000000000000000000000000000000010010000000000000; // D (0x0000000000012000) 
//    12'h77d : errs =          63'b000000000000000000000000000000000000000000000100010000000000000; // D (0x0000000000022000) 
//    12'h9fb : errs =          63'b000000000000000000000000000000000000000000001000010000000000000; // D (0x0000000000042000) 
//    12'h1ce : errs =          63'b000000000000000000000000000000000000000000010000010000000000000; // D (0x0000000000082000) 
//    12'h49d : errs =          63'b000000000000000000000000000000000000000000100000010000000000000; // D (0x0000000000102000) 
//    12'he3b : errs =          63'b000000000000000000000000000000000000000001000000010000000000000; // D (0x0000000000202000) 
//    12'he4e : errs =          63'b000000000000000000000000000000000000000010000000010000000000000; // D (0x0000000000402000) 
//    12'hea4 : errs =          63'b000000000000000000000000000000000000000100000000010000000000000; // D (0x0000000000802000) 
//    12'hf70 : errs =          63'b000000000000000000000000000000000000001000000000010000000000000; // D (0x0000000001002000) 
//    12'hcd8 : errs =          63'b000000000000000000000000000000000000010000000000010000000000000; // D (0x0000000002002000) 
//    12'hb88 : errs =          63'b000000000000000000000000000000000000100000000000010000000000000; // D (0x0000000004002000) 
//    12'h528 : errs =          63'b000000000000000000000000000000000001000000000000010000000000000; // D (0x0000000008002000) 
//    12'hd51 : errs =          63'b000000000000000000000000000000000010000000000000010000000000000; // D (0x0000000010002000) 
//    12'h89a : errs =          63'b000000000000000000000000000000000100000000000000010000000000000; // D (0x0000000020002000) 
//    12'h30c : errs =          63'b000000000000000000000000000000001000000000000000010000000000000; // D (0x0000000040002000) 
//    12'h119 : errs =          63'b000000000000000000000000000000010000000000000000010000000000000; // D (0x0000000080002000) 
//    12'h533 : errs =          63'b000000000000000000000000000000100000000000000000010000000000000; // D (0x0000000100002000) 
//    12'hd67 : errs =          63'b000000000000000000000000000001000000000000000000010000000000000; // D (0x0000000200002000) 
//    12'h8f6 : errs =          63'b000000000000000000000000000010000000000000000000010000000000000; // D (0x0000000400002000) 
//    12'h3d4 : errs =          63'b000000000000000000000000000100000000000000000000010000000000000; // D (0x0000000800002000) 
//    12'h0a9 : errs =          63'b000000000000000000000000001000000000000000000000010000000000000; // D (0x0000001000002000) 
//    12'h653 : errs =          63'b000000000000000000000000010000000000000000000000010000000000000; // D (0x0000002000002000) 
//    12'hba7 : errs =          63'b000000000000000000000000100000000000000000000000010000000000000; // D (0x0000004000002000) 
//    12'h576 : errs =          63'b000000000000000000000001000000000000000000000000010000000000000; // D (0x0000008000002000) 
//    12'hded : errs =          63'b000000000000000000000010000000000000000000000000010000000000000; // D (0x0000010000002000) 
//    12'h9e2 : errs =          63'b000000000000000000000100000000000000000000000000010000000000000; // D (0x0000020000002000) 
//    12'h1fc : errs =          63'b000000000000000000001000000000000000000000000000010000000000000; // D (0x0000040000002000) 
//    12'h4f9 : errs =          63'b000000000000000000010000000000000000000000000000010000000000000; // D (0x0000080000002000) 
//    12'hef3 : errs =          63'b000000000000000000100000000000000000000000000000010000000000000; // D (0x0000100000002000) 
//    12'hfde : errs =          63'b000000000000000001000000000000000000000000000000010000000000000; // D (0x0000200000002000) 
//    12'hd84 : errs =          63'b000000000000000010000000000000000000000000000000010000000000000; // D (0x0000400000002000) 
//    12'h930 : errs =          63'b000000000000000100000000000000000000000000000000010000000000000; // D (0x0000800000002000) 
//    12'h058 : errs =          63'b000000000000001000000000000000000000000000000000010000000000000; // D (0x0001000000002000) 
//    12'h7b1 : errs =          63'b000000000000010000000000000000000000000000000000010000000000000; // D (0x0002000000002000) 
//    12'h863 : errs =          63'b000000000000100000000000000000000000000000000000010000000000000; // D (0x0004000000002000) 
//    12'h2fe : errs =          63'b000000000001000000000000000000000000000000000000010000000000000; // D (0x0008000000002000) 
//    12'h2fd : errs =          63'b000000000010000000000000000000000000000000000000010000000000000; // D (0x0010000000002000) 
//    12'h2fb : errs =          63'b000000000100000000000000000000000000000000000000010000000000000; // D (0x0020000000002000) 
//    12'h2f7 : errs =          63'b000000001000000000000000000000000000000000000000010000000000000; // D (0x0040000000002000) 
//    12'h2ef : errs =          63'b000000010000000000000000000000000000000000000000010000000000000; // D (0x0080000000002000) 
//    12'h2df : errs =          63'b000000100000000000000000000000000000000000000000010000000000000; // D (0x0100000000002000) 
//    12'h2bf : errs =          63'b000001000000000000000000000000000000000000000000010000000000000; // D (0x0200000000002000) 
//    12'h27f : errs =          63'b000010000000000000000000000000000000000000000000010000000000000; // D (0x0400000000002000) 
//    12'h3ff : errs =          63'b000100000000000000000000000000000000000000000000010000000000000; // D (0x0800000000002000) 
//    12'h0ff : errs =          63'b001000000000000000000000000000000000000000000000010000000000000; // D (0x1000000000002000) 
//    12'h6ff : errs =          63'b010000000000000000000000000000000000000000000000010000000000000; // D (0x2000000000002000) 
//    12'haff : errs =          63'b100000000000000000000000000000000000000000000000010000000000000; // D (0x4000000000002000) 
    12'h0c7 : errs =          63'b000000000000000000000000000000000000000000000000100000000000001; // D (0x0000000000004001) 
    12'hf8c : errs =          63'b000000000000000000000000000000000000000000000000100000000000010; // D (0x0000000000004002) 
    12'h423 : errs =          63'b000000000000000000000000000000000000000000000000100000000000100; // D (0x0000000000004004) 
    12'h644 : errs =          63'b000000000000000000000000000000000000000000000000100000000001000; // D (0x0000000000004008) 
    12'h28a : errs =          63'b000000000000000000000000000000000000000000000000100000000010000; // D (0x0000000000004010) 
    12'hb16 : errs =          63'b000000000000000000000000000000000000000000000000100000000100000; // D (0x0000000000004020) 
    12'hd17 : errs =          63'b000000000000000000000000000000000000000000000000100000001000000; // D (0x0000000000004040) 
    12'h115 : errs =          63'b000000000000000000000000000000000000000000000000100000010000000; // D (0x0000000000004080) 
    12'hc28 : errs =          63'b000000000000000000000000000000000000000000000000100000100000000; // D (0x0000000000004100) 
    12'h36b : errs =          63'b000000000000000000000000000000000000000000000000100001000000000; // D (0x0000000000004200) 
    12'h8d4 : errs =          63'b000000000000000000000000000000000000000000000000100010000000000; // D (0x0000000000004400) 
    12'ha93 : errs =          63'b000000000000000000000000000000000000000000000000100100000000000; // D (0x0000000000004800) 
    12'he1d : errs =          63'b000000000000000000000000000000000000000000000000101000000000000; // D (0x0000000000005000) 
    12'h701 : errs =          63'b000000000000000000000000000000000000000000000000110000000000000; // D (0x0000000000006000) 
    12'h5fe : errs =          63'b000000000000000000000000000000000000000000000000100000000000000; // S (0x0000000000004000) 
//    12'he02 : errs =          63'b000000000000000000000000000000000000000000000001100000000000000; // D (0x000000000000c000) 
//    12'h73f : errs =          63'b000000000000000000000000000000000000000000000010100000000000000; // D (0x0000000000014000) 
//    12'h07c : errs =          63'b000000000000000000000000000000000000000000000100100000000000000; // D (0x0000000000024000) 
//    12'hefa : errs =          63'b000000000000000000000000000000000000000000001000100000000000000; // D (0x0000000000044000) 
//    12'h6cf : errs =          63'b000000000000000000000000000000000000000000010000100000000000000; // D (0x0000000000084000) 
//    12'h39c : errs =          63'b000000000000000000000000000000000000000000100000100000000000000; // D (0x0000000000104000) 
//    12'h93a : errs =          63'b000000000000000000000000000000000000000001000000100000000000000; // D (0x0000000000204000) 
//    12'h94f : errs =          63'b000000000000000000000000000000000000000010000000100000000000000; // D (0x0000000000404000) 
//    12'h9a5 : errs =          63'b000000000000000000000000000000000000000100000000100000000000000; // D (0x0000000000804000) 
//    12'h871 : errs =          63'b000000000000000000000000000000000000001000000000100000000000000; // D (0x0000000001004000) 
//    12'hbd9 : errs =          63'b000000000000000000000000000000000000010000000000100000000000000; // D (0x0000000002004000) 
//    12'hc89 : errs =          63'b000000000000000000000000000000000000100000000000100000000000000; // D (0x0000000004004000) 
//    12'h229 : errs =          63'b000000000000000000000000000000000001000000000000100000000000000; // D (0x0000000008004000) 
//    12'ha50 : errs =          63'b000000000000000000000000000000000010000000000000100000000000000; // D (0x0000000010004000) 
//    12'hf9b : errs =          63'b000000000000000000000000000000000100000000000000100000000000000; // D (0x0000000020004000) 
//    12'h40d : errs =          63'b000000000000000000000000000000001000000000000000100000000000000; // D (0x0000000040004000) 
//    12'h618 : errs =          63'b000000000000000000000000000000010000000000000000100000000000000; // D (0x0000000080004000) 
//    12'h232 : errs =          63'b000000000000000000000000000000100000000000000000100000000000000; // D (0x0000000100004000) 
//    12'ha66 : errs =          63'b000000000000000000000000000001000000000000000000100000000000000; // D (0x0000000200004000) 
//    12'hff7 : errs =          63'b000000000000000000000000000010000000000000000000100000000000000; // D (0x0000000400004000) 
//    12'h4d5 : errs =          63'b000000000000000000000000000100000000000000000000100000000000000; // D (0x0000000800004000) 
//    12'h7a8 : errs =          63'b000000000000000000000000001000000000000000000000100000000000000; // D (0x0000001000004000) 
//    12'h152 : errs =          63'b000000000000000000000000010000000000000000000000100000000000000; // D (0x0000002000004000) 
//    12'hca6 : errs =          63'b000000000000000000000000100000000000000000000000100000000000000; // D (0x0000004000004000) 
//    12'h277 : errs =          63'b000000000000000000000001000000000000000000000000100000000000000; // D (0x0000008000004000) 
//    12'haec : errs =          63'b000000000000000000000010000000000000000000000000100000000000000; // D (0x0000010000004000) 
//    12'hee3 : errs =          63'b000000000000000000000100000000000000000000000000100000000000000; // D (0x0000020000004000) 
//    12'h6fd : errs =          63'b000000000000000000001000000000000000000000000000100000000000000; // D (0x0000040000004000) 
//    12'h3f8 : errs =          63'b000000000000000000010000000000000000000000000000100000000000000; // D (0x0000080000004000) 
//    12'h9f2 : errs =          63'b000000000000000000100000000000000000000000000000100000000000000; // D (0x0000100000004000) 
//    12'h8df : errs =          63'b000000000000000001000000000000000000000000000000100000000000000; // D (0x0000200000004000) 
//    12'ha85 : errs =          63'b000000000000000010000000000000000000000000000000100000000000000; // D (0x0000400000004000) 
//    12'he31 : errs =          63'b000000000000000100000000000000000000000000000000100000000000000; // D (0x0000800000004000) 
//    12'h759 : errs =          63'b000000000000001000000000000000000000000000000000100000000000000; // D (0x0001000000004000) 
//    12'h0b0 : errs =          63'b000000000000010000000000000000000000000000000000100000000000000; // D (0x0002000000004000) 
//    12'hf62 : errs =          63'b000000000000100000000000000000000000000000000000100000000000000; // D (0x0004000000004000) 
//    12'h5ff : errs =          63'b000000000001000000000000000000000000000000000000100000000000000; // D (0x0008000000004000) 
//    12'h5fc : errs =          63'b000000000010000000000000000000000000000000000000100000000000000; // D (0x0010000000004000) 
//    12'h5fa : errs =          63'b000000000100000000000000000000000000000000000000100000000000000; // D (0x0020000000004000) 
//    12'h5f6 : errs =          63'b000000001000000000000000000000000000000000000000100000000000000; // D (0x0040000000004000) 
//    12'h5ee : errs =          63'b000000010000000000000000000000000000000000000000100000000000000; // D (0x0080000000004000) 
//    12'h5de : errs =          63'b000000100000000000000000000000000000000000000000100000000000000; // D (0x0100000000004000) 
//    12'h5be : errs =          63'b000001000000000000000000000000000000000000000000100000000000000; // D (0x0200000000004000) 
//    12'h57e : errs =          63'b000010000000000000000000000000000000000000000000100000000000000; // D (0x0400000000004000) 
//    12'h4fe : errs =          63'b000100000000000000000000000000000000000000000000100000000000000; // D (0x0800000000004000) 
//    12'h7fe : errs =          63'b001000000000000000000000000000000000000000000000100000000000000; // D (0x1000000000004000) 
//    12'h1fe : errs =          63'b010000000000000000000000000000000000000000000000100000000000000; // D (0x2000000000004000) 
//    12'hdfe : errs =          63'b100000000000000000000000000000000000000000000000100000000000000; // D (0x4000000000004000) 
    12'hec5 : errs =          63'b000000000000000000000000000000000000000000000001000000000000001; // D (0x0000000000008001) 
    12'h18e : errs =          63'b000000000000000000000000000000000000000000000001000000000000010; // D (0x0000000000008002) 
    12'ha21 : errs =          63'b000000000000000000000000000000000000000000000001000000000000100; // D (0x0000000000008004) 
    12'h846 : errs =          63'b000000000000000000000000000000000000000000000001000000000001000; // D (0x0000000000008008) 
    12'hc88 : errs =          63'b000000000000000000000000000000000000000000000001000000000010000; // D (0x0000000000008010) 
    12'h514 : errs =          63'b000000000000000000000000000000000000000000000001000000000100000; // D (0x0000000000008020) 
    12'h315 : errs =          63'b000000000000000000000000000000000000000000000001000000001000000; // D (0x0000000000008040) 
    12'hf17 : errs =          63'b000000000000000000000000000000000000000000000001000000010000000; // D (0x0000000000008080) 
    12'h22a : errs =          63'b000000000000000000000000000000000000000000000001000000100000000; // D (0x0000000000008100) 
    12'hd69 : errs =          63'b000000000000000000000000000000000000000000000001000001000000000; // D (0x0000000000008200) 
    12'h6d6 : errs =          63'b000000000000000000000000000000000000000000000001000010000000000; // D (0x0000000000008400) 
    12'h491 : errs =          63'b000000000000000000000000000000000000000000000001000100000000000; // D (0x0000000000008800) 
    12'h01f : errs =          63'b000000000000000000000000000000000000000000000001001000000000000; // D (0x0000000000009000) 
    12'h903 : errs =          63'b000000000000000000000000000000000000000000000001010000000000000; // D (0x000000000000a000) 
    12'he02 : errs =          63'b000000000000000000000000000000000000000000000001100000000000000; // D (0x000000000000c000) 
    12'hbfc : errs =          63'b000000000000000000000000000000000000000000000001000000000000000; // S (0x0000000000008000) 
//    12'h93d : errs =          63'b000000000000000000000000000000000000000000000011000000000000000; // D (0x0000000000018000) 
//    12'he7e : errs =          63'b000000000000000000000000000000000000000000000101000000000000000; // D (0x0000000000028000) 
//    12'h0f8 : errs =          63'b000000000000000000000000000000000000000000001001000000000000000; // D (0x0000000000048000) 
//    12'h8cd : errs =          63'b000000000000000000000000000000000000000000010001000000000000000; // D (0x0000000000088000) 
//    12'hd9e : errs =          63'b000000000000000000000000000000000000000000100001000000000000000; // D (0x0000000000108000) 
//    12'h738 : errs =          63'b000000000000000000000000000000000000000001000001000000000000000; // D (0x0000000000208000) 
//    12'h74d : errs =          63'b000000000000000000000000000000000000000010000001000000000000000; // D (0x0000000000408000) 
//    12'h7a7 : errs =          63'b000000000000000000000000000000000000000100000001000000000000000; // D (0x0000000000808000) 
//    12'h673 : errs =          63'b000000000000000000000000000000000000001000000001000000000000000; // D (0x0000000001008000) 
//    12'h5db : errs =          63'b000000000000000000000000000000000000010000000001000000000000000; // D (0x0000000002008000) 
//    12'h28b : errs =          63'b000000000000000000000000000000000000100000000001000000000000000; // D (0x0000000004008000) 
//    12'hc2b : errs =          63'b000000000000000000000000000000000001000000000001000000000000000; // D (0x0000000008008000) 
//    12'h452 : errs =          63'b000000000000000000000000000000000010000000000001000000000000000; // D (0x0000000010008000) 
//    12'h199 : errs =          63'b000000000000000000000000000000000100000000000001000000000000000; // D (0x0000000020008000) 
//    12'ha0f : errs =          63'b000000000000000000000000000000001000000000000001000000000000000; // D (0x0000000040008000) 
//    12'h81a : errs =          63'b000000000000000000000000000000010000000000000001000000000000000; // D (0x0000000080008000) 
//    12'hc30 : errs =          63'b000000000000000000000000000000100000000000000001000000000000000; // D (0x0000000100008000) 
//    12'h464 : errs =          63'b000000000000000000000000000001000000000000000001000000000000000; // D (0x0000000200008000) 
//    12'h1f5 : errs =          63'b000000000000000000000000000010000000000000000001000000000000000; // D (0x0000000400008000) 
//    12'had7 : errs =          63'b000000000000000000000000000100000000000000000001000000000000000; // D (0x0000000800008000) 
//    12'h9aa : errs =          63'b000000000000000000000000001000000000000000000001000000000000000; // D (0x0000001000008000) 
//    12'hf50 : errs =          63'b000000000000000000000000010000000000000000000001000000000000000; // D (0x0000002000008000) 
//    12'h2a4 : errs =          63'b000000000000000000000000100000000000000000000001000000000000000; // D (0x0000004000008000) 
//    12'hc75 : errs =          63'b000000000000000000000001000000000000000000000001000000000000000; // D (0x0000008000008000) 
//    12'h4ee : errs =          63'b000000000000000000000010000000000000000000000001000000000000000; // D (0x0000010000008000) 
//    12'h0e1 : errs =          63'b000000000000000000000100000000000000000000000001000000000000000; // D (0x0000020000008000) 
//    12'h8ff : errs =          63'b000000000000000000001000000000000000000000000001000000000000000; // D (0x0000040000008000) 
//    12'hdfa : errs =          63'b000000000000000000010000000000000000000000000001000000000000000; // D (0x0000080000008000) 
//    12'h7f0 : errs =          63'b000000000000000000100000000000000000000000000001000000000000000; // D (0x0000100000008000) 
//    12'h6dd : errs =          63'b000000000000000001000000000000000000000000000001000000000000000; // D (0x0000200000008000) 
//    12'h487 : errs =          63'b000000000000000010000000000000000000000000000001000000000000000; // D (0x0000400000008000) 
//    12'h033 : errs =          63'b000000000000000100000000000000000000000000000001000000000000000; // D (0x0000800000008000) 
//    12'h95b : errs =          63'b000000000000001000000000000000000000000000000001000000000000000; // D (0x0001000000008000) 
//    12'heb2 : errs =          63'b000000000000010000000000000000000000000000000001000000000000000; // D (0x0002000000008000) 
//    12'h160 : errs =          63'b000000000000100000000000000000000000000000000001000000000000000; // D (0x0004000000008000) 
//    12'hbfd : errs =          63'b000000000001000000000000000000000000000000000001000000000000000; // D (0x0008000000008000) 
//    12'hbfe : errs =          63'b000000000010000000000000000000000000000000000001000000000000000; // D (0x0010000000008000) 
//    12'hbf8 : errs =          63'b000000000100000000000000000000000000000000000001000000000000000; // D (0x0020000000008000) 
//    12'hbf4 : errs =          63'b000000001000000000000000000000000000000000000001000000000000000; // D (0x0040000000008000) 
//    12'hbec : errs =          63'b000000010000000000000000000000000000000000000001000000000000000; // D (0x0080000000008000) 
//    12'hbdc : errs =          63'b000000100000000000000000000000000000000000000001000000000000000; // D (0x0100000000008000) 
//    12'hbbc : errs =          63'b000001000000000000000000000000000000000000000001000000000000000; // D (0x0200000000008000) 
//    12'hb7c : errs =          63'b000010000000000000000000000000000000000000000001000000000000000; // D (0x0400000000008000) 
//    12'hafc : errs =          63'b000100000000000000000000000000000000000000000001000000000000000; // D (0x0800000000008000) 
//    12'h9fc : errs =          63'b001000000000000000000000000000000000000000000001000000000000000; // D (0x1000000000008000) 
//    12'hffc : errs =          63'b010000000000000000000000000000000000000000000001000000000000000; // D (0x2000000000008000) 
//    12'h3fc : errs =          63'b100000000000000000000000000000000000000000000001000000000000000; // D (0x4000000000008000) 
    12'h7f8 : errs =          63'b000000000000000000000000000000000000000000000010000000000000001; // D (0x0000000000010001) 
    12'h8b3 : errs =          63'b000000000000000000000000000000000000000000000010000000000000010; // D (0x0000000000010002) 
    12'h31c : errs =          63'b000000000000000000000000000000000000000000000010000000000000100; // D (0x0000000000010004) 
    12'h17b : errs =          63'b000000000000000000000000000000000000000000000010000000000001000; // D (0x0000000000010008) 
    12'h5b5 : errs =          63'b000000000000000000000000000000000000000000000010000000000010000; // D (0x0000000000010010) 
    12'hc29 : errs =          63'b000000000000000000000000000000000000000000000010000000000100000; // D (0x0000000000010020) 
    12'ha28 : errs =          63'b000000000000000000000000000000000000000000000010000000001000000; // D (0x0000000000010040) 
    12'h62a : errs =          63'b000000000000000000000000000000000000000000000010000000010000000; // D (0x0000000000010080) 
    12'hb17 : errs =          63'b000000000000000000000000000000000000000000000010000000100000000; // D (0x0000000000010100) 
    12'h454 : errs =          63'b000000000000000000000000000000000000000000000010000001000000000; // D (0x0000000000010200) 
    12'hfeb : errs =          63'b000000000000000000000000000000000000000000000010000010000000000; // D (0x0000000000010400) 
    12'hdac : errs =          63'b000000000000000000000000000000000000000000000010000100000000000; // D (0x0000000000010800) 
    12'h922 : errs =          63'b000000000000000000000000000000000000000000000010001000000000000; // D (0x0000000000011000) 
    12'h03e : errs =          63'b000000000000000000000000000000000000000000000010010000000000000; // D (0x0000000000012000) 
    12'h73f : errs =          63'b000000000000000000000000000000000000000000000010100000000000000; // D (0x0000000000014000) 
    12'h93d : errs =          63'b000000000000000000000000000000000000000000000011000000000000000; // D (0x0000000000018000) 
    12'h2c1 : errs =          63'b000000000000000000000000000000000000000000000010000000000000000; // S (0x0000000000010000) 
//    12'h743 : errs =          63'b000000000000000000000000000000000000000000000110000000000000000; // D (0x0000000000030000) 
//    12'h9c5 : errs =          63'b000000000000000000000000000000000000000000001010000000000000000; // D (0x0000000000050000) 
//    12'h1f0 : errs =          63'b000000000000000000000000000000000000000000010010000000000000000; // D (0x0000000000090000) 
//    12'h4a3 : errs =          63'b000000000000000000000000000000000000000000100010000000000000000; // D (0x0000000000110000) 
//    12'he05 : errs =          63'b000000000000000000000000000000000000000001000010000000000000000; // D (0x0000000000210000) 
//    12'he70 : errs =          63'b000000000000000000000000000000000000000010000010000000000000000; // D (0x0000000000410000) 
//    12'he9a : errs =          63'b000000000000000000000000000000000000000100000010000000000000000; // D (0x0000000000810000) 
//    12'hf4e : errs =          63'b000000000000000000000000000000000000001000000010000000000000000; // D (0x0000000001010000) 
//    12'hce6 : errs =          63'b000000000000000000000000000000000000010000000010000000000000000; // D (0x0000000002010000) 
//    12'hbb6 : errs =          63'b000000000000000000000000000000000000100000000010000000000000000; // D (0x0000000004010000) 
//    12'h516 : errs =          63'b000000000000000000000000000000000001000000000010000000000000000; // D (0x0000000008010000) 
//    12'hd6f : errs =          63'b000000000000000000000000000000000010000000000010000000000000000; // D (0x0000000010010000) 
//    12'h8a4 : errs =          63'b000000000000000000000000000000000100000000000010000000000000000; // D (0x0000000020010000) 
//    12'h332 : errs =          63'b000000000000000000000000000000001000000000000010000000000000000; // D (0x0000000040010000) 
//    12'h127 : errs =          63'b000000000000000000000000000000010000000000000010000000000000000; // D (0x0000000080010000) 
//    12'h50d : errs =          63'b000000000000000000000000000000100000000000000010000000000000000; // D (0x0000000100010000) 
//    12'hd59 : errs =          63'b000000000000000000000000000001000000000000000010000000000000000; // D (0x0000000200010000) 
//    12'h8c8 : errs =          63'b000000000000000000000000000010000000000000000010000000000000000; // D (0x0000000400010000) 
//    12'h3ea : errs =          63'b000000000000000000000000000100000000000000000010000000000000000; // D (0x0000000800010000) 
//    12'h097 : errs =          63'b000000000000000000000000001000000000000000000010000000000000000; // D (0x0000001000010000) 
//    12'h66d : errs =          63'b000000000000000000000000010000000000000000000010000000000000000; // D (0x0000002000010000) 
//    12'hb99 : errs =          63'b000000000000000000000000100000000000000000000010000000000000000; // D (0x0000004000010000) 
//    12'h548 : errs =          63'b000000000000000000000001000000000000000000000010000000000000000; // D (0x0000008000010000) 
//    12'hdd3 : errs =          63'b000000000000000000000010000000000000000000000010000000000000000; // D (0x0000010000010000) 
//    12'h9dc : errs =          63'b000000000000000000000100000000000000000000000010000000000000000; // D (0x0000020000010000) 
//    12'h1c2 : errs =          63'b000000000000000000001000000000000000000000000010000000000000000; // D (0x0000040000010000) 
//    12'h4c7 : errs =          63'b000000000000000000010000000000000000000000000010000000000000000; // D (0x0000080000010000) 
//    12'hecd : errs =          63'b000000000000000000100000000000000000000000000010000000000000000; // D (0x0000100000010000) 
//    12'hfe0 : errs =          63'b000000000000000001000000000000000000000000000010000000000000000; // D (0x0000200000010000) 
//    12'hdba : errs =          63'b000000000000000010000000000000000000000000000010000000000000000; // D (0x0000400000010000) 
//    12'h90e : errs =          63'b000000000000000100000000000000000000000000000010000000000000000; // D (0x0000800000010000) 
//    12'h066 : errs =          63'b000000000000001000000000000000000000000000000010000000000000000; // D (0x0001000000010000) 
//    12'h78f : errs =          63'b000000000000010000000000000000000000000000000010000000000000000; // D (0x0002000000010000) 
//    12'h85d : errs =          63'b000000000000100000000000000000000000000000000010000000000000000; // D (0x0004000000010000) 
//    12'h2c0 : errs =          63'b000000000001000000000000000000000000000000000010000000000000000; // D (0x0008000000010000) 
//    12'h2c3 : errs =          63'b000000000010000000000000000000000000000000000010000000000000000; // D (0x0010000000010000) 
//    12'h2c5 : errs =          63'b000000000100000000000000000000000000000000000010000000000000000; // D (0x0020000000010000) 
//    12'h2c9 : errs =          63'b000000001000000000000000000000000000000000000010000000000000000; // D (0x0040000000010000) 
//    12'h2d1 : errs =          63'b000000010000000000000000000000000000000000000010000000000000000; // D (0x0080000000010000) 
//    12'h2e1 : errs =          63'b000000100000000000000000000000000000000000000010000000000000000; // D (0x0100000000010000) 
//    12'h281 : errs =          63'b000001000000000000000000000000000000000000000010000000000000000; // D (0x0200000000010000) 
//    12'h241 : errs =          63'b000010000000000000000000000000000000000000000010000000000000000; // D (0x0400000000010000) 
//    12'h3c1 : errs =          63'b000100000000000000000000000000000000000000000010000000000000000; // D (0x0800000000010000) 
//    12'h0c1 : errs =          63'b001000000000000000000000000000000000000000000010000000000000000; // D (0x1000000000010000) 
//    12'h6c1 : errs =          63'b010000000000000000000000000000000000000000000010000000000000000; // D (0x2000000000010000) 
//    12'hac1 : errs =          63'b100000000000000000000000000000000000000000000010000000000000000; // D (0x4000000000010000) 
    12'h0bb : errs =          63'b000000000000000000000000000000000000000000000100000000000000001; // D (0x0000000000020001) 
    12'hff0 : errs =          63'b000000000000000000000000000000000000000000000100000000000000010; // D (0x0000000000020002) 
    12'h45f : errs =          63'b000000000000000000000000000000000000000000000100000000000000100; // D (0x0000000000020004) 
    12'h638 : errs =          63'b000000000000000000000000000000000000000000000100000000000001000; // D (0x0000000000020008) 
    12'h2f6 : errs =          63'b000000000000000000000000000000000000000000000100000000000010000; // D (0x0000000000020010) 
    12'hb6a : errs =          63'b000000000000000000000000000000000000000000000100000000000100000; // D (0x0000000000020020) 
    12'hd6b : errs =          63'b000000000000000000000000000000000000000000000100000000001000000; // D (0x0000000000020040) 
    12'h169 : errs =          63'b000000000000000000000000000000000000000000000100000000010000000; // D (0x0000000000020080) 
    12'hc54 : errs =          63'b000000000000000000000000000000000000000000000100000000100000000; // D (0x0000000000020100) 
    12'h317 : errs =          63'b000000000000000000000000000000000000000000000100000001000000000; // D (0x0000000000020200) 
    12'h8a8 : errs =          63'b000000000000000000000000000000000000000000000100000010000000000; // D (0x0000000000020400) 
    12'haef : errs =          63'b000000000000000000000000000000000000000000000100000100000000000; // D (0x0000000000020800) 
    12'he61 : errs =          63'b000000000000000000000000000000000000000000000100001000000000000; // D (0x0000000000021000) 
    12'h77d : errs =          63'b000000000000000000000000000000000000000000000100010000000000000; // D (0x0000000000022000) 
    12'h07c : errs =          63'b000000000000000000000000000000000000000000000100100000000000000; // D (0x0000000000024000) 
    12'he7e : errs =          63'b000000000000000000000000000000000000000000000101000000000000000; // D (0x0000000000028000) 
    12'h743 : errs =          63'b000000000000000000000000000000000000000000000110000000000000000; // D (0x0000000000030000) 
    12'h582 : errs =          63'b000000000000000000000000000000000000000000000100000000000000000; // S (0x0000000000020000) 
//    12'he86 : errs =          63'b000000000000000000000000000000000000000000001100000000000000000; // D (0x0000000000060000) 
//    12'h6b3 : errs =          63'b000000000000000000000000000000000000000000010100000000000000000; // D (0x00000000000a0000) 
//    12'h3e0 : errs =          63'b000000000000000000000000000000000000000000100100000000000000000; // D (0x0000000000120000) 
//    12'h946 : errs =          63'b000000000000000000000000000000000000000001000100000000000000000; // D (0x0000000000220000) 
//    12'h933 : errs =          63'b000000000000000000000000000000000000000010000100000000000000000; // D (0x0000000000420000) 
//    12'h9d9 : errs =          63'b000000000000000000000000000000000000000100000100000000000000000; // D (0x0000000000820000) 
//    12'h80d : errs =          63'b000000000000000000000000000000000000001000000100000000000000000; // D (0x0000000001020000) 
//    12'hba5 : errs =          63'b000000000000000000000000000000000000010000000100000000000000000; // D (0x0000000002020000) 
//    12'hcf5 : errs =          63'b000000000000000000000000000000000000100000000100000000000000000; // D (0x0000000004020000) 
//    12'h255 : errs =          63'b000000000000000000000000000000000001000000000100000000000000000; // D (0x0000000008020000) 
//    12'ha2c : errs =          63'b000000000000000000000000000000000010000000000100000000000000000; // D (0x0000000010020000) 
//    12'hfe7 : errs =          63'b000000000000000000000000000000000100000000000100000000000000000; // D (0x0000000020020000) 
//    12'h471 : errs =          63'b000000000000000000000000000000001000000000000100000000000000000; // D (0x0000000040020000) 
//    12'h664 : errs =          63'b000000000000000000000000000000010000000000000100000000000000000; // D (0x0000000080020000) 
//    12'h24e : errs =          63'b000000000000000000000000000000100000000000000100000000000000000; // D (0x0000000100020000) 
//    12'ha1a : errs =          63'b000000000000000000000000000001000000000000000100000000000000000; // D (0x0000000200020000) 
//    12'hf8b : errs =          63'b000000000000000000000000000010000000000000000100000000000000000; // D (0x0000000400020000) 
//    12'h4a9 : errs =          63'b000000000000000000000000000100000000000000000100000000000000000; // D (0x0000000800020000) 
//    12'h7d4 : errs =          63'b000000000000000000000000001000000000000000000100000000000000000; // D (0x0000001000020000) 
//    12'h12e : errs =          63'b000000000000000000000000010000000000000000000100000000000000000; // D (0x0000002000020000) 
//    12'hcda : errs =          63'b000000000000000000000000100000000000000000000100000000000000000; // D (0x0000004000020000) 
//    12'h20b : errs =          63'b000000000000000000000001000000000000000000000100000000000000000; // D (0x0000008000020000) 
//    12'ha90 : errs =          63'b000000000000000000000010000000000000000000000100000000000000000; // D (0x0000010000020000) 
//    12'he9f : errs =          63'b000000000000000000000100000000000000000000000100000000000000000; // D (0x0000020000020000) 
//    12'h681 : errs =          63'b000000000000000000001000000000000000000000000100000000000000000; // D (0x0000040000020000) 
//    12'h384 : errs =          63'b000000000000000000010000000000000000000000000100000000000000000; // D (0x0000080000020000) 
//    12'h98e : errs =          63'b000000000000000000100000000000000000000000000100000000000000000; // D (0x0000100000020000) 
//    12'h8a3 : errs =          63'b000000000000000001000000000000000000000000000100000000000000000; // D (0x0000200000020000) 
//    12'haf9 : errs =          63'b000000000000000010000000000000000000000000000100000000000000000; // D (0x0000400000020000) 
//    12'he4d : errs =          63'b000000000000000100000000000000000000000000000100000000000000000; // D (0x0000800000020000) 
//    12'h725 : errs =          63'b000000000000001000000000000000000000000000000100000000000000000; // D (0x0001000000020000) 
//    12'h0cc : errs =          63'b000000000000010000000000000000000000000000000100000000000000000; // D (0x0002000000020000) 
//    12'hf1e : errs =          63'b000000000000100000000000000000000000000000000100000000000000000; // D (0x0004000000020000) 
//    12'h583 : errs =          63'b000000000001000000000000000000000000000000000100000000000000000; // D (0x0008000000020000) 
//    12'h580 : errs =          63'b000000000010000000000000000000000000000000000100000000000000000; // D (0x0010000000020000) 
//    12'h586 : errs =          63'b000000000100000000000000000000000000000000000100000000000000000; // D (0x0020000000020000) 
//    12'h58a : errs =          63'b000000001000000000000000000000000000000000000100000000000000000; // D (0x0040000000020000) 
//    12'h592 : errs =          63'b000000010000000000000000000000000000000000000100000000000000000; // D (0x0080000000020000) 
//    12'h5a2 : errs =          63'b000000100000000000000000000000000000000000000100000000000000000; // D (0x0100000000020000) 
//    12'h5c2 : errs =          63'b000001000000000000000000000000000000000000000100000000000000000; // D (0x0200000000020000) 
//    12'h502 : errs =          63'b000010000000000000000000000000000000000000000100000000000000000; // D (0x0400000000020000) 
//    12'h482 : errs =          63'b000100000000000000000000000000000000000000000100000000000000000; // D (0x0800000000020000) 
//    12'h782 : errs =          63'b001000000000000000000000000000000000000000000100000000000000000; // D (0x1000000000020000) 
//    12'h182 : errs =          63'b010000000000000000000000000000000000000000000100000000000000000; // D (0x2000000000020000) 
//    12'hd82 : errs =          63'b100000000000000000000000000000000000000000000100000000000000000; // D (0x4000000000020000) 
    12'he3d : errs =          63'b000000000000000000000000000000000000000000001000000000000000001; // D (0x0000000000040001) 
    12'h176 : errs =          63'b000000000000000000000000000000000000000000001000000000000000010; // D (0x0000000000040002) 
    12'had9 : errs =          63'b000000000000000000000000000000000000000000001000000000000000100; // D (0x0000000000040004) 
    12'h8be : errs =          63'b000000000000000000000000000000000000000000001000000000000001000; // D (0x0000000000040008) 
    12'hc70 : errs =          63'b000000000000000000000000000000000000000000001000000000000010000; // D (0x0000000000040010) 
    12'h5ec : errs =          63'b000000000000000000000000000000000000000000001000000000000100000; // D (0x0000000000040020) 
    12'h3ed : errs =          63'b000000000000000000000000000000000000000000001000000000001000000; // D (0x0000000000040040) 
    12'hfef : errs =          63'b000000000000000000000000000000000000000000001000000000010000000; // D (0x0000000000040080) 
    12'h2d2 : errs =          63'b000000000000000000000000000000000000000000001000000000100000000; // D (0x0000000000040100) 
    12'hd91 : errs =          63'b000000000000000000000000000000000000000000001000000001000000000; // D (0x0000000000040200) 
    12'h62e : errs =          63'b000000000000000000000000000000000000000000001000000010000000000; // D (0x0000000000040400) 
    12'h469 : errs =          63'b000000000000000000000000000000000000000000001000000100000000000; // D (0x0000000000040800) 
    12'h0e7 : errs =          63'b000000000000000000000000000000000000000000001000001000000000000; // D (0x0000000000041000) 
    12'h9fb : errs =          63'b000000000000000000000000000000000000000000001000010000000000000; // D (0x0000000000042000) 
    12'hefa : errs =          63'b000000000000000000000000000000000000000000001000100000000000000; // D (0x0000000000044000) 
    12'h0f8 : errs =          63'b000000000000000000000000000000000000000000001001000000000000000; // D (0x0000000000048000) 
    12'h9c5 : errs =          63'b000000000000000000000000000000000000000000001010000000000000000; // D (0x0000000000050000) 
    12'he86 : errs =          63'b000000000000000000000000000000000000000000001100000000000000000; // D (0x0000000000060000) 
    12'hb04 : errs =          63'b000000000000000000000000000000000000000000001000000000000000000; // S (0x0000000000040000) 
//    12'h835 : errs =          63'b000000000000000000000000000000000000000000011000000000000000000; // D (0x00000000000c0000) 
//    12'hd66 : errs =          63'b000000000000000000000000000000000000000000101000000000000000000; // D (0x0000000000140000) 
//    12'h7c0 : errs =          63'b000000000000000000000000000000000000000001001000000000000000000; // D (0x0000000000240000) 
//    12'h7b5 : errs =          63'b000000000000000000000000000000000000000010001000000000000000000; // D (0x0000000000440000) 
//    12'h75f : errs =          63'b000000000000000000000000000000000000000100001000000000000000000; // D (0x0000000000840000) 
//    12'h68b : errs =          63'b000000000000000000000000000000000000001000001000000000000000000; // D (0x0000000001040000) 
//    12'h523 : errs =          63'b000000000000000000000000000000000000010000001000000000000000000; // D (0x0000000002040000) 
//    12'h273 : errs =          63'b000000000000000000000000000000000000100000001000000000000000000; // D (0x0000000004040000) 
//    12'hcd3 : errs =          63'b000000000000000000000000000000000001000000001000000000000000000; // D (0x0000000008040000) 
//    12'h4aa : errs =          63'b000000000000000000000000000000000010000000001000000000000000000; // D (0x0000000010040000) 
//    12'h161 : errs =          63'b000000000000000000000000000000000100000000001000000000000000000; // D (0x0000000020040000) 
//    12'haf7 : errs =          63'b000000000000000000000000000000001000000000001000000000000000000; // D (0x0000000040040000) 
//    12'h8e2 : errs =          63'b000000000000000000000000000000010000000000001000000000000000000; // D (0x0000000080040000) 
//    12'hcc8 : errs =          63'b000000000000000000000000000000100000000000001000000000000000000; // D (0x0000000100040000) 
//    12'h49c : errs =          63'b000000000000000000000000000001000000000000001000000000000000000; // D (0x0000000200040000) 
//    12'h10d : errs =          63'b000000000000000000000000000010000000000000001000000000000000000; // D (0x0000000400040000) 
//    12'ha2f : errs =          63'b000000000000000000000000000100000000000000001000000000000000000; // D (0x0000000800040000) 
//    12'h952 : errs =          63'b000000000000000000000000001000000000000000001000000000000000000; // D (0x0000001000040000) 
//    12'hfa8 : errs =          63'b000000000000000000000000010000000000000000001000000000000000000; // D (0x0000002000040000) 
//    12'h25c : errs =          63'b000000000000000000000000100000000000000000001000000000000000000; // D (0x0000004000040000) 
//    12'hc8d : errs =          63'b000000000000000000000001000000000000000000001000000000000000000; // D (0x0000008000040000) 
//    12'h416 : errs =          63'b000000000000000000000010000000000000000000001000000000000000000; // D (0x0000010000040000) 
//    12'h019 : errs =          63'b000000000000000000000100000000000000000000001000000000000000000; // D (0x0000020000040000) 
//    12'h807 : errs =          63'b000000000000000000001000000000000000000000001000000000000000000; // D (0x0000040000040000) 
//    12'hd02 : errs =          63'b000000000000000000010000000000000000000000001000000000000000000; // D (0x0000080000040000) 
//    12'h708 : errs =          63'b000000000000000000100000000000000000000000001000000000000000000; // D (0x0000100000040000) 
//    12'h625 : errs =          63'b000000000000000001000000000000000000000000001000000000000000000; // D (0x0000200000040000) 
//    12'h47f : errs =          63'b000000000000000010000000000000000000000000001000000000000000000; // D (0x0000400000040000) 
//    12'h0cb : errs =          63'b000000000000000100000000000000000000000000001000000000000000000; // D (0x0000800000040000) 
//    12'h9a3 : errs =          63'b000000000000001000000000000000000000000000001000000000000000000; // D (0x0001000000040000) 
//    12'he4a : errs =          63'b000000000000010000000000000000000000000000001000000000000000000; // D (0x0002000000040000) 
//    12'h198 : errs =          63'b000000000000100000000000000000000000000000001000000000000000000; // D (0x0004000000040000) 
//    12'hb05 : errs =          63'b000000000001000000000000000000000000000000001000000000000000000; // D (0x0008000000040000) 
//    12'hb06 : errs =          63'b000000000010000000000000000000000000000000001000000000000000000; // D (0x0010000000040000) 
//    12'hb00 : errs =          63'b000000000100000000000000000000000000000000001000000000000000000; // D (0x0020000000040000) 
//    12'hb0c : errs =          63'b000000001000000000000000000000000000000000001000000000000000000; // D (0x0040000000040000) 
//    12'hb14 : errs =          63'b000000010000000000000000000000000000000000001000000000000000000; // D (0x0080000000040000) 
//    12'hb24 : errs =          63'b000000100000000000000000000000000000000000001000000000000000000; // D (0x0100000000040000) 
//    12'hb44 : errs =          63'b000001000000000000000000000000000000000000001000000000000000000; // D (0x0200000000040000) 
//    12'hb84 : errs =          63'b000010000000000000000000000000000000000000001000000000000000000; // D (0x0400000000040000) 
//    12'ha04 : errs =          63'b000100000000000000000000000000000000000000001000000000000000000; // D (0x0800000000040000) 
//    12'h904 : errs =          63'b001000000000000000000000000000000000000000001000000000000000000; // D (0x1000000000040000) 
//    12'hf04 : errs =          63'b010000000000000000000000000000000000000000001000000000000000000; // D (0x2000000000040000) 
//    12'h304 : errs =          63'b100000000000000000000000000000000000000000001000000000000000000; // D (0x4000000000040000) 
    12'h608 : errs =          63'b000000000000000000000000000000000000000000010000000000000000001; // D (0x0000000000080001) 
    12'h943 : errs =          63'b000000000000000000000000000000000000000000010000000000000000010; // D (0x0000000000080002) 
    12'h2ec : errs =          63'b000000000000000000000000000000000000000000010000000000000000100; // D (0x0000000000080004) 
    12'h08b : errs =          63'b000000000000000000000000000000000000000000010000000000000001000; // D (0x0000000000080008) 
    12'h445 : errs =          63'b000000000000000000000000000000000000000000010000000000000010000; // D (0x0000000000080010) 
    12'hdd9 : errs =          63'b000000000000000000000000000000000000000000010000000000000100000; // D (0x0000000000080020) 
    12'hbd8 : errs =          63'b000000000000000000000000000000000000000000010000000000001000000; // D (0x0000000000080040) 
    12'h7da : errs =          63'b000000000000000000000000000000000000000000010000000000010000000; // D (0x0000000000080080) 
    12'hae7 : errs =          63'b000000000000000000000000000000000000000000010000000000100000000; // D (0x0000000000080100) 
    12'h5a4 : errs =          63'b000000000000000000000000000000000000000000010000000001000000000; // D (0x0000000000080200) 
    12'he1b : errs =          63'b000000000000000000000000000000000000000000010000000010000000000; // D (0x0000000000080400) 
    12'hc5c : errs =          63'b000000000000000000000000000000000000000000010000000100000000000; // D (0x0000000000080800) 
    12'h8d2 : errs =          63'b000000000000000000000000000000000000000000010000001000000000000; // D (0x0000000000081000) 
    12'h1ce : errs =          63'b000000000000000000000000000000000000000000010000010000000000000; // D (0x0000000000082000) 
    12'h6cf : errs =          63'b000000000000000000000000000000000000000000010000100000000000000; // D (0x0000000000084000) 
    12'h8cd : errs =          63'b000000000000000000000000000000000000000000010001000000000000000; // D (0x0000000000088000) 
    12'h1f0 : errs =          63'b000000000000000000000000000000000000000000010010000000000000000; // D (0x0000000000090000) 
    12'h6b3 : errs =          63'b000000000000000000000000000000000000000000010100000000000000000; // D (0x00000000000a0000) 
    12'h835 : errs =          63'b000000000000000000000000000000000000000000011000000000000000000; // D (0x00000000000c0000) 
    12'h331 : errs =          63'b000000000000000000000000000000000000000000010000000000000000000; // S (0x0000000000080000) 
//    12'h553 : errs =          63'b000000000000000000000000000000000000000000110000000000000000000; // D (0x0000000000180000) 
//    12'hff5 : errs =          63'b000000000000000000000000000000000000000001010000000000000000000; // D (0x0000000000280000) 
//    12'hf80 : errs =          63'b000000000000000000000000000000000000000010010000000000000000000; // D (0x0000000000480000) 
//    12'hf6a : errs =          63'b000000000000000000000000000000000000000100010000000000000000000; // D (0x0000000000880000) 
//    12'hebe : errs =          63'b000000000000000000000000000000000000001000010000000000000000000; // D (0x0000000001080000) 
//    12'hd16 : errs =          63'b000000000000000000000000000000000000010000010000000000000000000; // D (0x0000000002080000) 
//    12'ha46 : errs =          63'b000000000000000000000000000000000000100000010000000000000000000; // D (0x0000000004080000) 
//    12'h4e6 : errs =          63'b000000000000000000000000000000000001000000010000000000000000000; // D (0x0000000008080000) 
//    12'hc9f : errs =          63'b000000000000000000000000000000000010000000010000000000000000000; // D (0x0000000010080000) 
//    12'h954 : errs =          63'b000000000000000000000000000000000100000000010000000000000000000; // D (0x0000000020080000) 
//    12'h2c2 : errs =          63'b000000000000000000000000000000001000000000010000000000000000000; // D (0x0000000040080000) 
//    12'h0d7 : errs =          63'b000000000000000000000000000000010000000000010000000000000000000; // D (0x0000000080080000) 
//    12'h4fd : errs =          63'b000000000000000000000000000000100000000000010000000000000000000; // D (0x0000000100080000) 
//    12'hca9 : errs =          63'b000000000000000000000000000001000000000000010000000000000000000; // D (0x0000000200080000) 
//    12'h938 : errs =          63'b000000000000000000000000000010000000000000010000000000000000000; // D (0x0000000400080000) 
//    12'h21a : errs =          63'b000000000000000000000000000100000000000000010000000000000000000; // D (0x0000000800080000) 
//    12'h167 : errs =          63'b000000000000000000000000001000000000000000010000000000000000000; // D (0x0000001000080000) 
//    12'h79d : errs =          63'b000000000000000000000000010000000000000000010000000000000000000; // D (0x0000002000080000) 
//    12'ha69 : errs =          63'b000000000000000000000000100000000000000000010000000000000000000; // D (0x0000004000080000) 
//    12'h4b8 : errs =          63'b000000000000000000000001000000000000000000010000000000000000000; // D (0x0000008000080000) 
//    12'hc23 : errs =          63'b000000000000000000000010000000000000000000010000000000000000000; // D (0x0000010000080000) 
//    12'h82c : errs =          63'b000000000000000000000100000000000000000000010000000000000000000; // D (0x0000020000080000) 
//    12'h032 : errs =          63'b000000000000000000001000000000000000000000010000000000000000000; // D (0x0000040000080000) 
//    12'h537 : errs =          63'b000000000000000000010000000000000000000000010000000000000000000; // D (0x0000080000080000) 
//    12'hf3d : errs =          63'b000000000000000000100000000000000000000000010000000000000000000; // D (0x0000100000080000) 
//    12'he10 : errs =          63'b000000000000000001000000000000000000000000010000000000000000000; // D (0x0000200000080000) 
//    12'hc4a : errs =          63'b000000000000000010000000000000000000000000010000000000000000000; // D (0x0000400000080000) 
//    12'h8fe : errs =          63'b000000000000000100000000000000000000000000010000000000000000000; // D (0x0000800000080000) 
//    12'h196 : errs =          63'b000000000000001000000000000000000000000000010000000000000000000; // D (0x0001000000080000) 
//    12'h67f : errs =          63'b000000000000010000000000000000000000000000010000000000000000000; // D (0x0002000000080000) 
//    12'h9ad : errs =          63'b000000000000100000000000000000000000000000010000000000000000000; // D (0x0004000000080000) 
//    12'h330 : errs =          63'b000000000001000000000000000000000000000000010000000000000000000; // D (0x0008000000080000) 
//    12'h333 : errs =          63'b000000000010000000000000000000000000000000010000000000000000000; // D (0x0010000000080000) 
//    12'h335 : errs =          63'b000000000100000000000000000000000000000000010000000000000000000; // D (0x0020000000080000) 
//    12'h339 : errs =          63'b000000001000000000000000000000000000000000010000000000000000000; // D (0x0040000000080000) 
//    12'h321 : errs =          63'b000000010000000000000000000000000000000000010000000000000000000; // D (0x0080000000080000) 
//    12'h311 : errs =          63'b000000100000000000000000000000000000000000010000000000000000000; // D (0x0100000000080000) 
//    12'h371 : errs =          63'b000001000000000000000000000000000000000000010000000000000000000; // D (0x0200000000080000) 
//    12'h3b1 : errs =          63'b000010000000000000000000000000000000000000010000000000000000000; // D (0x0400000000080000) 
//    12'h231 : errs =          63'b000100000000000000000000000000000000000000010000000000000000000; // D (0x0800000000080000) 
//    12'h131 : errs =          63'b001000000000000000000000000000000000000000010000000000000000000; // D (0x1000000000080000) 
//    12'h731 : errs =          63'b010000000000000000000000000000000000000000010000000000000000000; // D (0x2000000000080000) 
//    12'hb31 : errs =          63'b100000000000000000000000000000000000000000010000000000000000000; // D (0x4000000000080000) 
    12'h35b : errs =          63'b000000000000000000000000000000000000000000100000000000000000001; // D (0x0000000000100001) 
    12'hc10 : errs =          63'b000000000000000000000000000000000000000000100000000000000000010; // D (0x0000000000100002) 
    12'h7bf : errs =          63'b000000000000000000000000000000000000000000100000000000000000100; // D (0x0000000000100004) 
    12'h5d8 : errs =          63'b000000000000000000000000000000000000000000100000000000000001000; // D (0x0000000000100008) 
    12'h116 : errs =          63'b000000000000000000000000000000000000000000100000000000000010000; // D (0x0000000000100010) 
    12'h88a : errs =          63'b000000000000000000000000000000000000000000100000000000000100000; // D (0x0000000000100020) 
    12'he8b : errs =          63'b000000000000000000000000000000000000000000100000000000001000000; // D (0x0000000000100040) 
    12'h289 : errs =          63'b000000000000000000000000000000000000000000100000000000010000000; // D (0x0000000000100080) 
    12'hfb4 : errs =          63'b000000000000000000000000000000000000000000100000000000100000000; // D (0x0000000000100100) 
    12'h0f7 : errs =          63'b000000000000000000000000000000000000000000100000000001000000000; // D (0x0000000000100200) 
    12'hb48 : errs =          63'b000000000000000000000000000000000000000000100000000010000000000; // D (0x0000000000100400) 
    12'h90f : errs =          63'b000000000000000000000000000000000000000000100000000100000000000; // D (0x0000000000100800) 
    12'hd81 : errs =          63'b000000000000000000000000000000000000000000100000001000000000000; // D (0x0000000000101000) 
    12'h49d : errs =          63'b000000000000000000000000000000000000000000100000010000000000000; // D (0x0000000000102000) 
    12'h39c : errs =          63'b000000000000000000000000000000000000000000100000100000000000000; // D (0x0000000000104000) 
    12'hd9e : errs =          63'b000000000000000000000000000000000000000000100001000000000000000; // D (0x0000000000108000) 
    12'h4a3 : errs =          63'b000000000000000000000000000000000000000000100010000000000000000; // D (0x0000000000110000) 
    12'h3e0 : errs =          63'b000000000000000000000000000000000000000000100100000000000000000; // D (0x0000000000120000) 
    12'hd66 : errs =          63'b000000000000000000000000000000000000000000101000000000000000000; // D (0x0000000000140000) 
    12'h553 : errs =          63'b000000000000000000000000000000000000000000110000000000000000000; // D (0x0000000000180000) 
    12'h662 : errs =          63'b000000000000000000000000000000000000000000100000000000000000000; // S (0x0000000000100000) 
//    12'haa6 : errs =          63'b000000000000000000000000000000000000000001100000000000000000000; // D (0x0000000000300000) 
//    12'had3 : errs =          63'b000000000000000000000000000000000000000010100000000000000000000; // D (0x0000000000500000) 
//    12'ha39 : errs =          63'b000000000000000000000000000000000000000100100000000000000000000; // D (0x0000000000900000) 
//    12'hbed : errs =          63'b000000000000000000000000000000000000001000100000000000000000000; // D (0x0000000001100000) 
//    12'h845 : errs =          63'b000000000000000000000000000000000000010000100000000000000000000; // D (0x0000000002100000) 
//    12'hf15 : errs =          63'b000000000000000000000000000000000000100000100000000000000000000; // D (0x0000000004100000) 
//    12'h1b5 : errs =          63'b000000000000000000000000000000000001000000100000000000000000000; // D (0x0000000008100000) 
//    12'h9cc : errs =          63'b000000000000000000000000000000000010000000100000000000000000000; // D (0x0000000010100000) 
//    12'hc07 : errs =          63'b000000000000000000000000000000000100000000100000000000000000000; // D (0x0000000020100000) 
//    12'h791 : errs =          63'b000000000000000000000000000000001000000000100000000000000000000; // D (0x0000000040100000) 
//    12'h584 : errs =          63'b000000000000000000000000000000010000000000100000000000000000000; // D (0x0000000080100000) 
//    12'h1ae : errs =          63'b000000000000000000000000000000100000000000100000000000000000000; // D (0x0000000100100000) 
//    12'h9fa : errs =          63'b000000000000000000000000000001000000000000100000000000000000000; // D (0x0000000200100000) 
//    12'hc6b : errs =          63'b000000000000000000000000000010000000000000100000000000000000000; // D (0x0000000400100000) 
//    12'h749 : errs =          63'b000000000000000000000000000100000000000000100000000000000000000; // D (0x0000000800100000) 
//    12'h434 : errs =          63'b000000000000000000000000001000000000000000100000000000000000000; // D (0x0000001000100000) 
//    12'h2ce : errs =          63'b000000000000000000000000010000000000000000100000000000000000000; // D (0x0000002000100000) 
//    12'hf3a : errs =          63'b000000000000000000000000100000000000000000100000000000000000000; // D (0x0000004000100000) 
//    12'h1eb : errs =          63'b000000000000000000000001000000000000000000100000000000000000000; // D (0x0000008000100000) 
//    12'h970 : errs =          63'b000000000000000000000010000000000000000000100000000000000000000; // D (0x0000010000100000) 
//    12'hd7f : errs =          63'b000000000000000000000100000000000000000000100000000000000000000; // D (0x0000020000100000) 
//    12'h561 : errs =          63'b000000000000000000001000000000000000000000100000000000000000000; // D (0x0000040000100000) 
//    12'h064 : errs =          63'b000000000000000000010000000000000000000000100000000000000000000; // D (0x0000080000100000) 
//    12'ha6e : errs =          63'b000000000000000000100000000000000000000000100000000000000000000; // D (0x0000100000100000) 
//    12'hb43 : errs =          63'b000000000000000001000000000000000000000000100000000000000000000; // D (0x0000200000100000) 
//    12'h919 : errs =          63'b000000000000000010000000000000000000000000100000000000000000000; // D (0x0000400000100000) 
//    12'hdad : errs =          63'b000000000000000100000000000000000000000000100000000000000000000; // D (0x0000800000100000) 
//    12'h4c5 : errs =          63'b000000000000001000000000000000000000000000100000000000000000000; // D (0x0001000000100000) 
//    12'h32c : errs =          63'b000000000000010000000000000000000000000000100000000000000000000; // D (0x0002000000100000) 
//    12'hcfe : errs =          63'b000000000000100000000000000000000000000000100000000000000000000; // D (0x0004000000100000) 
//    12'h663 : errs =          63'b000000000001000000000000000000000000000000100000000000000000000; // D (0x0008000000100000) 
//    12'h660 : errs =          63'b000000000010000000000000000000000000000000100000000000000000000; // D (0x0010000000100000) 
//    12'h666 : errs =          63'b000000000100000000000000000000000000000000100000000000000000000; // D (0x0020000000100000) 
//    12'h66a : errs =          63'b000000001000000000000000000000000000000000100000000000000000000; // D (0x0040000000100000) 
//    12'h672 : errs =          63'b000000010000000000000000000000000000000000100000000000000000000; // D (0x0080000000100000) 
//    12'h642 : errs =          63'b000000100000000000000000000000000000000000100000000000000000000; // D (0x0100000000100000) 
//    12'h622 : errs =          63'b000001000000000000000000000000000000000000100000000000000000000; // D (0x0200000000100000) 
//    12'h6e2 : errs =          63'b000010000000000000000000000000000000000000100000000000000000000; // D (0x0400000000100000) 
//    12'h762 : errs =          63'b000100000000000000000000000000000000000000100000000000000000000; // D (0x0800000000100000) 
//    12'h462 : errs =          63'b001000000000000000000000000000000000000000100000000000000000000; // D (0x1000000000100000) 
//    12'h262 : errs =          63'b010000000000000000000000000000000000000000100000000000000000000; // D (0x2000000000100000) 
//    12'he62 : errs =          63'b100000000000000000000000000000000000000000100000000000000000000; // D (0x4000000000100000) 
    12'h9fd : errs =          63'b000000000000000000000000000000000000000001000000000000000000001; // D (0x0000000000200001) 
    12'h6b6 : errs =          63'b000000000000000000000000000000000000000001000000000000000000010; // D (0x0000000000200002) 
    12'hd19 : errs =          63'b000000000000000000000000000000000000000001000000000000000000100; // D (0x0000000000200004) 
    12'hf7e : errs =          63'b000000000000000000000000000000000000000001000000000000000001000; // D (0x0000000000200008) 
    12'hbb0 : errs =          63'b000000000000000000000000000000000000000001000000000000000010000; // D (0x0000000000200010) 
    12'h22c : errs =          63'b000000000000000000000000000000000000000001000000000000000100000; // D (0x0000000000200020) 
    12'h42d : errs =          63'b000000000000000000000000000000000000000001000000000000001000000; // D (0x0000000000200040) 
    12'h82f : errs =          63'b000000000000000000000000000000000000000001000000000000010000000; // D (0x0000000000200080) 
    12'h512 : errs =          63'b000000000000000000000000000000000000000001000000000000100000000; // D (0x0000000000200100) 
    12'ha51 : errs =          63'b000000000000000000000000000000000000000001000000000001000000000; // D (0x0000000000200200) 
    12'h1ee : errs =          63'b000000000000000000000000000000000000000001000000000010000000000; // D (0x0000000000200400) 
    12'h3a9 : errs =          63'b000000000000000000000000000000000000000001000000000100000000000; // D (0x0000000000200800) 
    12'h727 : errs =          63'b000000000000000000000000000000000000000001000000001000000000000; // D (0x0000000000201000) 
    12'he3b : errs =          63'b000000000000000000000000000000000000000001000000010000000000000; // D (0x0000000000202000) 
    12'h93a : errs =          63'b000000000000000000000000000000000000000001000000100000000000000; // D (0x0000000000204000) 
    12'h738 : errs =          63'b000000000000000000000000000000000000000001000001000000000000000; // D (0x0000000000208000) 
    12'he05 : errs =          63'b000000000000000000000000000000000000000001000010000000000000000; // D (0x0000000000210000) 
    12'h946 : errs =          63'b000000000000000000000000000000000000000001000100000000000000000; // D (0x0000000000220000) 
    12'h7c0 : errs =          63'b000000000000000000000000000000000000000001001000000000000000000; // D (0x0000000000240000) 
    12'hff5 : errs =          63'b000000000000000000000000000000000000000001010000000000000000000; // D (0x0000000000280000) 
    12'haa6 : errs =          63'b000000000000000000000000000000000000000001100000000000000000000; // D (0x0000000000300000) 
    12'hcc4 : errs =          63'b000000000000000000000000000000000000000001000000000000000000000; // S (0x0000000000200000) 
//    12'h075 : errs =          63'b000000000000000000000000000000000000000011000000000000000000000; // D (0x0000000000600000) 
//    12'h09f : errs =          63'b000000000000000000000000000000000000000101000000000000000000000; // D (0x0000000000a00000) 
//    12'h14b : errs =          63'b000000000000000000000000000000000000001001000000000000000000000; // D (0x0000000001200000) 
//    12'h2e3 : errs =          63'b000000000000000000000000000000000000010001000000000000000000000; // D (0x0000000002200000) 
//    12'h5b3 : errs =          63'b000000000000000000000000000000000000100001000000000000000000000; // D (0x0000000004200000) 
//    12'hb13 : errs =          63'b000000000000000000000000000000000001000001000000000000000000000; // D (0x0000000008200000) 
//    12'h36a : errs =          63'b000000000000000000000000000000000010000001000000000000000000000; // D (0x0000000010200000) 
//    12'h6a1 : errs =          63'b000000000000000000000000000000000100000001000000000000000000000; // D (0x0000000020200000) 
//    12'hd37 : errs =          63'b000000000000000000000000000000001000000001000000000000000000000; // D (0x0000000040200000) 
//    12'hf22 : errs =          63'b000000000000000000000000000000010000000001000000000000000000000; // D (0x0000000080200000) 
//    12'hb08 : errs =          63'b000000000000000000000000000000100000000001000000000000000000000; // D (0x0000000100200000) 
//    12'h35c : errs =          63'b000000000000000000000000000001000000000001000000000000000000000; // D (0x0000000200200000) 
//    12'h6cd : errs =          63'b000000000000000000000000000010000000000001000000000000000000000; // D (0x0000000400200000) 
//    12'hdef : errs =          63'b000000000000000000000000000100000000000001000000000000000000000; // D (0x0000000800200000) 
//    12'he92 : errs =          63'b000000000000000000000000001000000000000001000000000000000000000; // D (0x0000001000200000) 
//    12'h868 : errs =          63'b000000000000000000000000010000000000000001000000000000000000000; // D (0x0000002000200000) 
//    12'h59c : errs =          63'b000000000000000000000000100000000000000001000000000000000000000; // D (0x0000004000200000) 
//    12'hb4d : errs =          63'b000000000000000000000001000000000000000001000000000000000000000; // D (0x0000008000200000) 
//    12'h3d6 : errs =          63'b000000000000000000000010000000000000000001000000000000000000000; // D (0x0000010000200000) 
//    12'h7d9 : errs =          63'b000000000000000000000100000000000000000001000000000000000000000; // D (0x0000020000200000) 
//    12'hfc7 : errs =          63'b000000000000000000001000000000000000000001000000000000000000000; // D (0x0000040000200000) 
//    12'hac2 : errs =          63'b000000000000000000010000000000000000000001000000000000000000000; // D (0x0000080000200000) 
//    12'h0c8 : errs =          63'b000000000000000000100000000000000000000001000000000000000000000; // D (0x0000100000200000) 
//    12'h1e5 : errs =          63'b000000000000000001000000000000000000000001000000000000000000000; // D (0x0000200000200000) 
//    12'h3bf : errs =          63'b000000000000000010000000000000000000000001000000000000000000000; // D (0x0000400000200000) 
//    12'h70b : errs =          63'b000000000000000100000000000000000000000001000000000000000000000; // D (0x0000800000200000) 
//    12'he63 : errs =          63'b000000000000001000000000000000000000000001000000000000000000000; // D (0x0001000000200000) 
//    12'h98a : errs =          63'b000000000000010000000000000000000000000001000000000000000000000; // D (0x0002000000200000) 
//    12'h658 : errs =          63'b000000000000100000000000000000000000000001000000000000000000000; // D (0x0004000000200000) 
//    12'hcc5 : errs =          63'b000000000001000000000000000000000000000001000000000000000000000; // D (0x0008000000200000) 
//    12'hcc6 : errs =          63'b000000000010000000000000000000000000000001000000000000000000000; // D (0x0010000000200000) 
//    12'hcc0 : errs =          63'b000000000100000000000000000000000000000001000000000000000000000; // D (0x0020000000200000) 
//    12'hccc : errs =          63'b000000001000000000000000000000000000000001000000000000000000000; // D (0x0040000000200000) 
//    12'hcd4 : errs =          63'b000000010000000000000000000000000000000001000000000000000000000; // D (0x0080000000200000) 
//    12'hce4 : errs =          63'b000000100000000000000000000000000000000001000000000000000000000; // D (0x0100000000200000) 
//    12'hc84 : errs =          63'b000001000000000000000000000000000000000001000000000000000000000; // D (0x0200000000200000) 
//    12'hc44 : errs =          63'b000010000000000000000000000000000000000001000000000000000000000; // D (0x0400000000200000) 
//    12'hdc4 : errs =          63'b000100000000000000000000000000000000000001000000000000000000000; // D (0x0800000000200000) 
//    12'hec4 : errs =          63'b001000000000000000000000000000000000000001000000000000000000000; // D (0x1000000000200000) 
//    12'h8c4 : errs =          63'b010000000000000000000000000000000000000001000000000000000000000; // D (0x2000000000200000) 
//    12'h4c4 : errs =          63'b100000000000000000000000000000000000000001000000000000000000000; // D (0x4000000000200000) 
    12'h988 : errs =          63'b000000000000000000000000000000000000000010000000000000000000001; // D (0x0000000000400001) 
    12'h6c3 : errs =          63'b000000000000000000000000000000000000000010000000000000000000010; // D (0x0000000000400002) 
    12'hd6c : errs =          63'b000000000000000000000000000000000000000010000000000000000000100; // D (0x0000000000400004) 
    12'hf0b : errs =          63'b000000000000000000000000000000000000000010000000000000000001000; // D (0x0000000000400008) 
    12'hbc5 : errs =          63'b000000000000000000000000000000000000000010000000000000000010000; // D (0x0000000000400010) 
    12'h259 : errs =          63'b000000000000000000000000000000000000000010000000000000000100000; // D (0x0000000000400020) 
    12'h458 : errs =          63'b000000000000000000000000000000000000000010000000000000001000000; // D (0x0000000000400040) 
    12'h85a : errs =          63'b000000000000000000000000000000000000000010000000000000010000000; // D (0x0000000000400080) 
    12'h567 : errs =          63'b000000000000000000000000000000000000000010000000000000100000000; // D (0x0000000000400100) 
    12'ha24 : errs =          63'b000000000000000000000000000000000000000010000000000001000000000; // D (0x0000000000400200) 
    12'h19b : errs =          63'b000000000000000000000000000000000000000010000000000010000000000; // D (0x0000000000400400) 
    12'h3dc : errs =          63'b000000000000000000000000000000000000000010000000000100000000000; // D (0x0000000000400800) 
    12'h752 : errs =          63'b000000000000000000000000000000000000000010000000001000000000000; // D (0x0000000000401000) 
    12'he4e : errs =          63'b000000000000000000000000000000000000000010000000010000000000000; // D (0x0000000000402000) 
    12'h94f : errs =          63'b000000000000000000000000000000000000000010000000100000000000000; // D (0x0000000000404000) 
    12'h74d : errs =          63'b000000000000000000000000000000000000000010000001000000000000000; // D (0x0000000000408000) 
    12'he70 : errs =          63'b000000000000000000000000000000000000000010000010000000000000000; // D (0x0000000000410000) 
    12'h933 : errs =          63'b000000000000000000000000000000000000000010000100000000000000000; // D (0x0000000000420000) 
    12'h7b5 : errs =          63'b000000000000000000000000000000000000000010001000000000000000000; // D (0x0000000000440000) 
    12'hf80 : errs =          63'b000000000000000000000000000000000000000010010000000000000000000; // D (0x0000000000480000) 
    12'had3 : errs =          63'b000000000000000000000000000000000000000010100000000000000000000; // D (0x0000000000500000) 
    12'h075 : errs =          63'b000000000000000000000000000000000000000011000000000000000000000; // D (0x0000000000600000) 
    12'hcb1 : errs =          63'b000000000000000000000000000000000000000010000000000000000000000; // S (0x0000000000400000) 
//    12'h0ea : errs =          63'b000000000000000000000000000000000000000110000000000000000000000; // D (0x0000000000c00000) 
//    12'h13e : errs =          63'b000000000000000000000000000000000000001010000000000000000000000; // D (0x0000000001400000) 
//    12'h296 : errs =          63'b000000000000000000000000000000000000010010000000000000000000000; // D (0x0000000002400000) 
//    12'h5c6 : errs =          63'b000000000000000000000000000000000000100010000000000000000000000; // D (0x0000000004400000) 
//    12'hb66 : errs =          63'b000000000000000000000000000000000001000010000000000000000000000; // D (0x0000000008400000) 
//    12'h31f : errs =          63'b000000000000000000000000000000000010000010000000000000000000000; // D (0x0000000010400000) 
//    12'h6d4 : errs =          63'b000000000000000000000000000000000100000010000000000000000000000; // D (0x0000000020400000) 
//    12'hd42 : errs =          63'b000000000000000000000000000000001000000010000000000000000000000; // D (0x0000000040400000) 
//    12'hf57 : errs =          63'b000000000000000000000000000000010000000010000000000000000000000; // D (0x0000000080400000) 
//    12'hb7d : errs =          63'b000000000000000000000000000000100000000010000000000000000000000; // D (0x0000000100400000) 
//    12'h329 : errs =          63'b000000000000000000000000000001000000000010000000000000000000000; // D (0x0000000200400000) 
//    12'h6b8 : errs =          63'b000000000000000000000000000010000000000010000000000000000000000; // D (0x0000000400400000) 
//    12'hd9a : errs =          63'b000000000000000000000000000100000000000010000000000000000000000; // D (0x0000000800400000) 
//    12'hee7 : errs =          63'b000000000000000000000000001000000000000010000000000000000000000; // D (0x0000001000400000) 
//    12'h81d : errs =          63'b000000000000000000000000010000000000000010000000000000000000000; // D (0x0000002000400000) 
//    12'h5e9 : errs =          63'b000000000000000000000000100000000000000010000000000000000000000; // D (0x0000004000400000) 
//    12'hb38 : errs =          63'b000000000000000000000001000000000000000010000000000000000000000; // D (0x0000008000400000) 
//    12'h3a3 : errs =          63'b000000000000000000000010000000000000000010000000000000000000000; // D (0x0000010000400000) 
//    12'h7ac : errs =          63'b000000000000000000000100000000000000000010000000000000000000000; // D (0x0000020000400000) 
//    12'hfb2 : errs =          63'b000000000000000000001000000000000000000010000000000000000000000; // D (0x0000040000400000) 
//    12'hab7 : errs =          63'b000000000000000000010000000000000000000010000000000000000000000; // D (0x0000080000400000) 
//    12'h0bd : errs =          63'b000000000000000000100000000000000000000010000000000000000000000; // D (0x0000100000400000) 
//    12'h190 : errs =          63'b000000000000000001000000000000000000000010000000000000000000000; // D (0x0000200000400000) 
//    12'h3ca : errs =          63'b000000000000000010000000000000000000000010000000000000000000000; // D (0x0000400000400000) 
//    12'h77e : errs =          63'b000000000000000100000000000000000000000010000000000000000000000; // D (0x0000800000400000) 
//    12'he16 : errs =          63'b000000000000001000000000000000000000000010000000000000000000000; // D (0x0001000000400000) 
//    12'h9ff : errs =          63'b000000000000010000000000000000000000000010000000000000000000000; // D (0x0002000000400000) 
//    12'h62d : errs =          63'b000000000000100000000000000000000000000010000000000000000000000; // D (0x0004000000400000) 
//    12'hcb0 : errs =          63'b000000000001000000000000000000000000000010000000000000000000000; // D (0x0008000000400000) 
//    12'hcb3 : errs =          63'b000000000010000000000000000000000000000010000000000000000000000; // D (0x0010000000400000) 
//    12'hcb5 : errs =          63'b000000000100000000000000000000000000000010000000000000000000000; // D (0x0020000000400000) 
//    12'hcb9 : errs =          63'b000000001000000000000000000000000000000010000000000000000000000; // D (0x0040000000400000) 
//    12'hca1 : errs =          63'b000000010000000000000000000000000000000010000000000000000000000; // D (0x0080000000400000) 
//    12'hc91 : errs =          63'b000000100000000000000000000000000000000010000000000000000000000; // D (0x0100000000400000) 
//    12'hcf1 : errs =          63'b000001000000000000000000000000000000000010000000000000000000000; // D (0x0200000000400000) 
//    12'hc31 : errs =          63'b000010000000000000000000000000000000000010000000000000000000000; // D (0x0400000000400000) 
//    12'hdb1 : errs =          63'b000100000000000000000000000000000000000010000000000000000000000; // D (0x0800000000400000) 
//    12'heb1 : errs =          63'b001000000000000000000000000000000000000010000000000000000000000; // D (0x1000000000400000) 
//    12'h8b1 : errs =          63'b010000000000000000000000000000000000000010000000000000000000000; // D (0x2000000000400000) 
//    12'h4b1 : errs =          63'b100000000000000000000000000000000000000010000000000000000000000; // D (0x4000000000400000) 
    12'h962 : errs =          63'b000000000000000000000000000000000000000100000000000000000000001; // D (0x0000000000800001) 
    12'h629 : errs =          63'b000000000000000000000000000000000000000100000000000000000000010; // D (0x0000000000800002) 
    12'hd86 : errs =          63'b000000000000000000000000000000000000000100000000000000000000100; // D (0x0000000000800004) 
    12'hfe1 : errs =          63'b000000000000000000000000000000000000000100000000000000000001000; // D (0x0000000000800008) 
    12'hb2f : errs =          63'b000000000000000000000000000000000000000100000000000000000010000; // D (0x0000000000800010) 
    12'h2b3 : errs =          63'b000000000000000000000000000000000000000100000000000000000100000; // D (0x0000000000800020) 
    12'h4b2 : errs =          63'b000000000000000000000000000000000000000100000000000000001000000; // D (0x0000000000800040) 
    12'h8b0 : errs =          63'b000000000000000000000000000000000000000100000000000000010000000; // D (0x0000000000800080) 
    12'h58d : errs =          63'b000000000000000000000000000000000000000100000000000000100000000; // D (0x0000000000800100) 
    12'hace : errs =          63'b000000000000000000000000000000000000000100000000000001000000000; // D (0x0000000000800200) 
    12'h171 : errs =          63'b000000000000000000000000000000000000000100000000000010000000000; // D (0x0000000000800400) 
    12'h336 : errs =          63'b000000000000000000000000000000000000000100000000000100000000000; // D (0x0000000000800800) 
    12'h7b8 : errs =          63'b000000000000000000000000000000000000000100000000001000000000000; // D (0x0000000000801000) 
    12'hea4 : errs =          63'b000000000000000000000000000000000000000100000000010000000000000; // D (0x0000000000802000) 
    12'h9a5 : errs =          63'b000000000000000000000000000000000000000100000000100000000000000; // D (0x0000000000804000) 
    12'h7a7 : errs =          63'b000000000000000000000000000000000000000100000001000000000000000; // D (0x0000000000808000) 
    12'he9a : errs =          63'b000000000000000000000000000000000000000100000010000000000000000; // D (0x0000000000810000) 
    12'h9d9 : errs =          63'b000000000000000000000000000000000000000100000100000000000000000; // D (0x0000000000820000) 
    12'h75f : errs =          63'b000000000000000000000000000000000000000100001000000000000000000; // D (0x0000000000840000) 
    12'hf6a : errs =          63'b000000000000000000000000000000000000000100010000000000000000000; // D (0x0000000000880000) 
    12'ha39 : errs =          63'b000000000000000000000000000000000000000100100000000000000000000; // D (0x0000000000900000) 
    12'h09f : errs =          63'b000000000000000000000000000000000000000101000000000000000000000; // D (0x0000000000a00000) 
    12'h0ea : errs =          63'b000000000000000000000000000000000000000110000000000000000000000; // D (0x0000000000c00000) 
    12'hc5b : errs =          63'b000000000000000000000000000000000000000100000000000000000000000; // S (0x0000000000800000) 
//    12'h1d4 : errs =          63'b000000000000000000000000000000000000001100000000000000000000000; // D (0x0000000001800000) 
//    12'h27c : errs =          63'b000000000000000000000000000000000000010100000000000000000000000; // D (0x0000000002800000) 
//    12'h52c : errs =          63'b000000000000000000000000000000000000100100000000000000000000000; // D (0x0000000004800000) 
//    12'hb8c : errs =          63'b000000000000000000000000000000000001000100000000000000000000000; // D (0x0000000008800000) 
//    12'h3f5 : errs =          63'b000000000000000000000000000000000010000100000000000000000000000; // D (0x0000000010800000) 
//    12'h63e : errs =          63'b000000000000000000000000000000000100000100000000000000000000000; // D (0x0000000020800000) 
//    12'hda8 : errs =          63'b000000000000000000000000000000001000000100000000000000000000000; // D (0x0000000040800000) 
//    12'hfbd : errs =          63'b000000000000000000000000000000010000000100000000000000000000000; // D (0x0000000080800000) 
//    12'hb97 : errs =          63'b000000000000000000000000000000100000000100000000000000000000000; // D (0x0000000100800000) 
//    12'h3c3 : errs =          63'b000000000000000000000000000001000000000100000000000000000000000; // D (0x0000000200800000) 
//    12'h652 : errs =          63'b000000000000000000000000000010000000000100000000000000000000000; // D (0x0000000400800000) 
//    12'hd70 : errs =          63'b000000000000000000000000000100000000000100000000000000000000000; // D (0x0000000800800000) 
//    12'he0d : errs =          63'b000000000000000000000000001000000000000100000000000000000000000; // D (0x0000001000800000) 
//    12'h8f7 : errs =          63'b000000000000000000000000010000000000000100000000000000000000000; // D (0x0000002000800000) 
//    12'h503 : errs =          63'b000000000000000000000000100000000000000100000000000000000000000; // D (0x0000004000800000) 
//    12'hbd2 : errs =          63'b000000000000000000000001000000000000000100000000000000000000000; // D (0x0000008000800000) 
//    12'h349 : errs =          63'b000000000000000000000010000000000000000100000000000000000000000; // D (0x0000010000800000) 
//    12'h746 : errs =          63'b000000000000000000000100000000000000000100000000000000000000000; // D (0x0000020000800000) 
//    12'hf58 : errs =          63'b000000000000000000001000000000000000000100000000000000000000000; // D (0x0000040000800000) 
//    12'ha5d : errs =          63'b000000000000000000010000000000000000000100000000000000000000000; // D (0x0000080000800000) 
//    12'h057 : errs =          63'b000000000000000000100000000000000000000100000000000000000000000; // D (0x0000100000800000) 
//    12'h17a : errs =          63'b000000000000000001000000000000000000000100000000000000000000000; // D (0x0000200000800000) 
//    12'h320 : errs =          63'b000000000000000010000000000000000000000100000000000000000000000; // D (0x0000400000800000) 
//    12'h794 : errs =          63'b000000000000000100000000000000000000000100000000000000000000000; // D (0x0000800000800000) 
//    12'hefc : errs =          63'b000000000000001000000000000000000000000100000000000000000000000; // D (0x0001000000800000) 
//    12'h915 : errs =          63'b000000000000010000000000000000000000000100000000000000000000000; // D (0x0002000000800000) 
//    12'h6c7 : errs =          63'b000000000000100000000000000000000000000100000000000000000000000; // D (0x0004000000800000) 
//    12'hc5a : errs =          63'b000000000001000000000000000000000000000100000000000000000000000; // D (0x0008000000800000) 
//    12'hc59 : errs =          63'b000000000010000000000000000000000000000100000000000000000000000; // D (0x0010000000800000) 
//    12'hc5f : errs =          63'b000000000100000000000000000000000000000100000000000000000000000; // D (0x0020000000800000) 
//    12'hc53 : errs =          63'b000000001000000000000000000000000000000100000000000000000000000; // D (0x0040000000800000) 
//    12'hc4b : errs =          63'b000000010000000000000000000000000000000100000000000000000000000; // D (0x0080000000800000) 
//    12'hc7b : errs =          63'b000000100000000000000000000000000000000100000000000000000000000; // D (0x0100000000800000) 
//    12'hc1b : errs =          63'b000001000000000000000000000000000000000100000000000000000000000; // D (0x0200000000800000) 
//    12'hcdb : errs =          63'b000010000000000000000000000000000000000100000000000000000000000; // D (0x0400000000800000) 
//    12'hd5b : errs =          63'b000100000000000000000000000000000000000100000000000000000000000; // D (0x0800000000800000) 
//    12'he5b : errs =          63'b001000000000000000000000000000000000000100000000000000000000000; // D (0x1000000000800000) 
//    12'h85b : errs =          63'b010000000000000000000000000000000000000100000000000000000000000; // D (0x2000000000800000) 
//    12'h45b : errs =          63'b100000000000000000000000000000000000000100000000000000000000000; // D (0x4000000000800000) 
    12'h8b6 : errs =          63'b000000000000000000000000000000000000001000000000000000000000001; // D (0x0000000001000001) 
    12'h7fd : errs =          63'b000000000000000000000000000000000000001000000000000000000000010; // D (0x0000000001000002) 
    12'hc52 : errs =          63'b000000000000000000000000000000000000001000000000000000000000100; // D (0x0000000001000004) 
    12'he35 : errs =          63'b000000000000000000000000000000000000001000000000000000000001000; // D (0x0000000001000008) 
    12'hafb : errs =          63'b000000000000000000000000000000000000001000000000000000000010000; // D (0x0000000001000010) 
    12'h367 : errs =          63'b000000000000000000000000000000000000001000000000000000000100000; // D (0x0000000001000020) 
    12'h566 : errs =          63'b000000000000000000000000000000000000001000000000000000001000000; // D (0x0000000001000040) 
    12'h964 : errs =          63'b000000000000000000000000000000000000001000000000000000010000000; // D (0x0000000001000080) 
    12'h459 : errs =          63'b000000000000000000000000000000000000001000000000000000100000000; // D (0x0000000001000100) 
    12'hb1a : errs =          63'b000000000000000000000000000000000000001000000000000001000000000; // D (0x0000000001000200) 
    12'h0a5 : errs =          63'b000000000000000000000000000000000000001000000000000010000000000; // D (0x0000000001000400) 
    12'h2e2 : errs =          63'b000000000000000000000000000000000000001000000000000100000000000; // D (0x0000000001000800) 
    12'h66c : errs =          63'b000000000000000000000000000000000000001000000000001000000000000; // D (0x0000000001001000) 
    12'hf70 : errs =          63'b000000000000000000000000000000000000001000000000010000000000000; // D (0x0000000001002000) 
    12'h871 : errs =          63'b000000000000000000000000000000000000001000000000100000000000000; // D (0x0000000001004000) 
    12'h673 : errs =          63'b000000000000000000000000000000000000001000000001000000000000000; // D (0x0000000001008000) 
    12'hf4e : errs =          63'b000000000000000000000000000000000000001000000010000000000000000; // D (0x0000000001010000) 
    12'h80d : errs =          63'b000000000000000000000000000000000000001000000100000000000000000; // D (0x0000000001020000) 
    12'h68b : errs =          63'b000000000000000000000000000000000000001000001000000000000000000; // D (0x0000000001040000) 
    12'hebe : errs =          63'b000000000000000000000000000000000000001000010000000000000000000; // D (0x0000000001080000) 
    12'hbed : errs =          63'b000000000000000000000000000000000000001000100000000000000000000; // D (0x0000000001100000) 
    12'h14b : errs =          63'b000000000000000000000000000000000000001001000000000000000000000; // D (0x0000000001200000) 
    12'h13e : errs =          63'b000000000000000000000000000000000000001010000000000000000000000; // D (0x0000000001400000) 
    12'h1d4 : errs =          63'b000000000000000000000000000000000000001100000000000000000000000; // D (0x0000000001800000) 
    12'hd8f : errs =          63'b000000000000000000000000000000000000001000000000000000000000000; // S (0x0000000001000000) 
//    12'h3a8 : errs =          63'b000000000000000000000000000000000000011000000000000000000000000; // D (0x0000000003000000) 
//    12'h4f8 : errs =          63'b000000000000000000000000000000000000101000000000000000000000000; // D (0x0000000005000000) 
//    12'ha58 : errs =          63'b000000000000000000000000000000000001001000000000000000000000000; // D (0x0000000009000000) 
//    12'h221 : errs =          63'b000000000000000000000000000000000010001000000000000000000000000; // D (0x0000000011000000) 
//    12'h7ea : errs =          63'b000000000000000000000000000000000100001000000000000000000000000; // D (0x0000000021000000) 
//    12'hc7c : errs =          63'b000000000000000000000000000000001000001000000000000000000000000; // D (0x0000000041000000) 
//    12'he69 : errs =          63'b000000000000000000000000000000010000001000000000000000000000000; // D (0x0000000081000000) 
//    12'ha43 : errs =          63'b000000000000000000000000000000100000001000000000000000000000000; // D (0x0000000101000000) 
//    12'h217 : errs =          63'b000000000000000000000000000001000000001000000000000000000000000; // D (0x0000000201000000) 
//    12'h786 : errs =          63'b000000000000000000000000000010000000001000000000000000000000000; // D (0x0000000401000000) 
//    12'hca4 : errs =          63'b000000000000000000000000000100000000001000000000000000000000000; // D (0x0000000801000000) 
//    12'hfd9 : errs =          63'b000000000000000000000000001000000000001000000000000000000000000; // D (0x0000001001000000) 
//    12'h923 : errs =          63'b000000000000000000000000010000000000001000000000000000000000000; // D (0x0000002001000000) 
//    12'h4d7 : errs =          63'b000000000000000000000000100000000000001000000000000000000000000; // D (0x0000004001000000) 
//    12'ha06 : errs =          63'b000000000000000000000001000000000000001000000000000000000000000; // D (0x0000008001000000) 
//    12'h29d : errs =          63'b000000000000000000000010000000000000001000000000000000000000000; // D (0x0000010001000000) 
//    12'h692 : errs =          63'b000000000000000000000100000000000000001000000000000000000000000; // D (0x0000020001000000) 
//    12'he8c : errs =          63'b000000000000000000001000000000000000001000000000000000000000000; // D (0x0000040001000000) 
//    12'hb89 : errs =          63'b000000000000000000010000000000000000001000000000000000000000000; // D (0x0000080001000000) 
//    12'h183 : errs =          63'b000000000000000000100000000000000000001000000000000000000000000; // D (0x0000100001000000) 
//    12'h0ae : errs =          63'b000000000000000001000000000000000000001000000000000000000000000; // D (0x0000200001000000) 
//    12'h2f4 : errs =          63'b000000000000000010000000000000000000001000000000000000000000000; // D (0x0000400001000000) 
//    12'h640 : errs =          63'b000000000000000100000000000000000000001000000000000000000000000; // D (0x0000800001000000) 
//    12'hf28 : errs =          63'b000000000000001000000000000000000000001000000000000000000000000; // D (0x0001000001000000) 
//    12'h8c1 : errs =          63'b000000000000010000000000000000000000001000000000000000000000000; // D (0x0002000001000000) 
//    12'h713 : errs =          63'b000000000000100000000000000000000000001000000000000000000000000; // D (0x0004000001000000) 
//    12'hd8e : errs =          63'b000000000001000000000000000000000000001000000000000000000000000; // D (0x0008000001000000) 
//    12'hd8d : errs =          63'b000000000010000000000000000000000000001000000000000000000000000; // D (0x0010000001000000) 
//    12'hd8b : errs =          63'b000000000100000000000000000000000000001000000000000000000000000; // D (0x0020000001000000) 
//    12'hd87 : errs =          63'b000000001000000000000000000000000000001000000000000000000000000; // D (0x0040000001000000) 
//    12'hd9f : errs =          63'b000000010000000000000000000000000000001000000000000000000000000; // D (0x0080000001000000) 
//    12'hdaf : errs =          63'b000000100000000000000000000000000000001000000000000000000000000; // D (0x0100000001000000) 
//    12'hdcf : errs =          63'b000001000000000000000000000000000000001000000000000000000000000; // D (0x0200000001000000) 
//    12'hd0f : errs =          63'b000010000000000000000000000000000000001000000000000000000000000; // D (0x0400000001000000) 
//    12'hc8f : errs =          63'b000100000000000000000000000000000000001000000000000000000000000; // D (0x0800000001000000) 
//    12'hf8f : errs =          63'b001000000000000000000000000000000000001000000000000000000000000; // D (0x1000000001000000) 
//    12'h98f : errs =          63'b010000000000000000000000000000000000001000000000000000000000000; // D (0x2000000001000000) 
//    12'h58f : errs =          63'b100000000000000000000000000000000000001000000000000000000000000; // D (0x4000000001000000) 
    12'hb1e : errs =          63'b000000000000000000000000000000000000010000000000000000000000001; // D (0x0000000002000001) 
    12'h455 : errs =          63'b000000000000000000000000000000000000010000000000000000000000010; // D (0x0000000002000002) 
    12'hffa : errs =          63'b000000000000000000000000000000000000010000000000000000000000100; // D (0x0000000002000004) 
    12'hd9d : errs =          63'b000000000000000000000000000000000000010000000000000000000001000; // D (0x0000000002000008) 
    12'h953 : errs =          63'b000000000000000000000000000000000000010000000000000000000010000; // D (0x0000000002000010) 
    12'h0cf : errs =          63'b000000000000000000000000000000000000010000000000000000000100000; // D (0x0000000002000020) 
    12'h6ce : errs =          63'b000000000000000000000000000000000000010000000000000000001000000; // D (0x0000000002000040) 
    12'hacc : errs =          63'b000000000000000000000000000000000000010000000000000000010000000; // D (0x0000000002000080) 
    12'h7f1 : errs =          63'b000000000000000000000000000000000000010000000000000000100000000; // D (0x0000000002000100) 
    12'h8b2 : errs =          63'b000000000000000000000000000000000000010000000000000001000000000; // D (0x0000000002000200) 
    12'h30d : errs =          63'b000000000000000000000000000000000000010000000000000010000000000; // D (0x0000000002000400) 
    12'h14a : errs =          63'b000000000000000000000000000000000000010000000000000100000000000; // D (0x0000000002000800) 
    12'h5c4 : errs =          63'b000000000000000000000000000000000000010000000000001000000000000; // D (0x0000000002001000) 
    12'hcd8 : errs =          63'b000000000000000000000000000000000000010000000000010000000000000; // D (0x0000000002002000) 
    12'hbd9 : errs =          63'b000000000000000000000000000000000000010000000000100000000000000; // D (0x0000000002004000) 
    12'h5db : errs =          63'b000000000000000000000000000000000000010000000001000000000000000; // D (0x0000000002008000) 
    12'hce6 : errs =          63'b000000000000000000000000000000000000010000000010000000000000000; // D (0x0000000002010000) 
    12'hba5 : errs =          63'b000000000000000000000000000000000000010000000100000000000000000; // D (0x0000000002020000) 
    12'h523 : errs =          63'b000000000000000000000000000000000000010000001000000000000000000; // D (0x0000000002040000) 
    12'hd16 : errs =          63'b000000000000000000000000000000000000010000010000000000000000000; // D (0x0000000002080000) 
    12'h845 : errs =          63'b000000000000000000000000000000000000010000100000000000000000000; // D (0x0000000002100000) 
    12'h2e3 : errs =          63'b000000000000000000000000000000000000010001000000000000000000000; // D (0x0000000002200000) 
    12'h296 : errs =          63'b000000000000000000000000000000000000010010000000000000000000000; // D (0x0000000002400000) 
    12'h27c : errs =          63'b000000000000000000000000000000000000010100000000000000000000000; // D (0x0000000002800000) 
    12'h3a8 : errs =          63'b000000000000000000000000000000000000011000000000000000000000000; // D (0x0000000003000000) 
    12'he27 : errs =          63'b000000000000000000000000000000000000010000000000000000000000000; // S (0x0000000002000000) 
//    12'h750 : errs =          63'b000000000000000000000000000000000000110000000000000000000000000; // D (0x0000000006000000) 
//    12'h9f0 : errs =          63'b000000000000000000000000000000000001010000000000000000000000000; // D (0x000000000a000000) 
//    12'h189 : errs =          63'b000000000000000000000000000000000010010000000000000000000000000; // D (0x0000000012000000) 
//    12'h442 : errs =          63'b000000000000000000000000000000000100010000000000000000000000000; // D (0x0000000022000000) 
//    12'hfd4 : errs =          63'b000000000000000000000000000000001000010000000000000000000000000; // D (0x0000000042000000) 
//    12'hdc1 : errs =          63'b000000000000000000000000000000010000010000000000000000000000000; // D (0x0000000082000000) 
//    12'h9eb : errs =          63'b000000000000000000000000000000100000010000000000000000000000000; // D (0x0000000102000000) 
//    12'h1bf : errs =          63'b000000000000000000000000000001000000010000000000000000000000000; // D (0x0000000202000000) 
//    12'h42e : errs =          63'b000000000000000000000000000010000000010000000000000000000000000; // D (0x0000000402000000) 
//    12'hf0c : errs =          63'b000000000000000000000000000100000000010000000000000000000000000; // D (0x0000000802000000) 
//    12'hc71 : errs =          63'b000000000000000000000000001000000000010000000000000000000000000; // D (0x0000001002000000) 
//    12'ha8b : errs =          63'b000000000000000000000000010000000000010000000000000000000000000; // D (0x0000002002000000) 
//    12'h77f : errs =          63'b000000000000000000000000100000000000010000000000000000000000000; // D (0x0000004002000000) 
//    12'h9ae : errs =          63'b000000000000000000000001000000000000010000000000000000000000000; // D (0x0000008002000000) 
//    12'h135 : errs =          63'b000000000000000000000010000000000000010000000000000000000000000; // D (0x0000010002000000) 
//    12'h53a : errs =          63'b000000000000000000000100000000000000010000000000000000000000000; // D (0x0000020002000000) 
//    12'hd24 : errs =          63'b000000000000000000001000000000000000010000000000000000000000000; // D (0x0000040002000000) 
//    12'h821 : errs =          63'b000000000000000000010000000000000000010000000000000000000000000; // D (0x0000080002000000) 
//    12'h22b : errs =          63'b000000000000000000100000000000000000010000000000000000000000000; // D (0x0000100002000000) 
//    12'h306 : errs =          63'b000000000000000001000000000000000000010000000000000000000000000; // D (0x0000200002000000) 
//    12'h15c : errs =          63'b000000000000000010000000000000000000010000000000000000000000000; // D (0x0000400002000000) 
//    12'h5e8 : errs =          63'b000000000000000100000000000000000000010000000000000000000000000; // D (0x0000800002000000) 
//    12'hc80 : errs =          63'b000000000000001000000000000000000000010000000000000000000000000; // D (0x0001000002000000) 
//    12'hb69 : errs =          63'b000000000000010000000000000000000000010000000000000000000000000; // D (0x0002000002000000) 
//    12'h4bb : errs =          63'b000000000000100000000000000000000000010000000000000000000000000; // D (0x0004000002000000) 
//    12'he26 : errs =          63'b000000000001000000000000000000000000010000000000000000000000000; // D (0x0008000002000000) 
//    12'he25 : errs =          63'b000000000010000000000000000000000000010000000000000000000000000; // D (0x0010000002000000) 
//    12'he23 : errs =          63'b000000000100000000000000000000000000010000000000000000000000000; // D (0x0020000002000000) 
//    12'he2f : errs =          63'b000000001000000000000000000000000000010000000000000000000000000; // D (0x0040000002000000) 
//    12'he37 : errs =          63'b000000010000000000000000000000000000010000000000000000000000000; // D (0x0080000002000000) 
//    12'he07 : errs =          63'b000000100000000000000000000000000000010000000000000000000000000; // D (0x0100000002000000) 
//    12'he67 : errs =          63'b000001000000000000000000000000000000010000000000000000000000000; // D (0x0200000002000000) 
//    12'hea7 : errs =          63'b000010000000000000000000000000000000010000000000000000000000000; // D (0x0400000002000000) 
//    12'hf27 : errs =          63'b000100000000000000000000000000000000010000000000000000000000000; // D (0x0800000002000000) 
//    12'hc27 : errs =          63'b001000000000000000000000000000000000010000000000000000000000000; // D (0x1000000002000000) 
//    12'ha27 : errs =          63'b010000000000000000000000000000000000010000000000000000000000000; // D (0x2000000002000000) 
//    12'h627 : errs =          63'b100000000000000000000000000000000000010000000000000000000000000; // D (0x4000000002000000) 
    12'hc4e : errs =          63'b000000000000000000000000000000000000100000000000000000000000001; // D (0x0000000004000001) 
    12'h305 : errs =          63'b000000000000000000000000000000000000100000000000000000000000010; // D (0x0000000004000002) 
    12'h8aa : errs =          63'b000000000000000000000000000000000000100000000000000000000000100; // D (0x0000000004000004) 
    12'hacd : errs =          63'b000000000000000000000000000000000000100000000000000000000001000; // D (0x0000000004000008) 
    12'he03 : errs =          63'b000000000000000000000000000000000000100000000000000000000010000; // D (0x0000000004000010) 
    12'h79f : errs =          63'b000000000000000000000000000000000000100000000000000000000100000; // D (0x0000000004000020) 
    12'h19e : errs =          63'b000000000000000000000000000000000000100000000000000000001000000; // D (0x0000000004000040) 
    12'hd9c : errs =          63'b000000000000000000000000000000000000100000000000000000010000000; // D (0x0000000004000080) 
    12'h0a1 : errs =          63'b000000000000000000000000000000000000100000000000000000100000000; // D (0x0000000004000100) 
    12'hfe2 : errs =          63'b000000000000000000000000000000000000100000000000000001000000000; // D (0x0000000004000200) 
    12'h45d : errs =          63'b000000000000000000000000000000000000100000000000000010000000000; // D (0x0000000004000400) 
    12'h61a : errs =          63'b000000000000000000000000000000000000100000000000000100000000000; // D (0x0000000004000800) 
    12'h294 : errs =          63'b000000000000000000000000000000000000100000000000001000000000000; // D (0x0000000004001000) 
    12'hb88 : errs =          63'b000000000000000000000000000000000000100000000000010000000000000; // D (0x0000000004002000) 
    12'hc89 : errs =          63'b000000000000000000000000000000000000100000000000100000000000000; // D (0x0000000004004000) 
    12'h28b : errs =          63'b000000000000000000000000000000000000100000000001000000000000000; // D (0x0000000004008000) 
    12'hbb6 : errs =          63'b000000000000000000000000000000000000100000000010000000000000000; // D (0x0000000004010000) 
    12'hcf5 : errs =          63'b000000000000000000000000000000000000100000000100000000000000000; // D (0x0000000004020000) 
    12'h273 : errs =          63'b000000000000000000000000000000000000100000001000000000000000000; // D (0x0000000004040000) 
    12'ha46 : errs =          63'b000000000000000000000000000000000000100000010000000000000000000; // D (0x0000000004080000) 
    12'hf15 : errs =          63'b000000000000000000000000000000000000100000100000000000000000000; // D (0x0000000004100000) 
    12'h5b3 : errs =          63'b000000000000000000000000000000000000100001000000000000000000000; // D (0x0000000004200000) 
    12'h5c6 : errs =          63'b000000000000000000000000000000000000100010000000000000000000000; // D (0x0000000004400000) 
    12'h52c : errs =          63'b000000000000000000000000000000000000100100000000000000000000000; // D (0x0000000004800000) 
    12'h4f8 : errs =          63'b000000000000000000000000000000000000101000000000000000000000000; // D (0x0000000005000000) 
    12'h750 : errs =          63'b000000000000000000000000000000000000110000000000000000000000000; // D (0x0000000006000000) 
    12'h977 : errs =          63'b000000000000000000000000000000000000100000000000000000000000000; // S (0x0000000004000000) 
//    12'hea0 : errs =          63'b000000000000000000000000000000000001100000000000000000000000000; // D (0x000000000c000000) 
//    12'h6d9 : errs =          63'b000000000000000000000000000000000010100000000000000000000000000; // D (0x0000000014000000) 
//    12'h312 : errs =          63'b000000000000000000000000000000000100100000000000000000000000000; // D (0x0000000024000000) 
//    12'h884 : errs =          63'b000000000000000000000000000000001000100000000000000000000000000; // D (0x0000000044000000) 
//    12'ha91 : errs =          63'b000000000000000000000000000000010000100000000000000000000000000; // D (0x0000000084000000) 
//    12'hebb : errs =          63'b000000000000000000000000000000100000100000000000000000000000000; // D (0x0000000104000000) 
//    12'h6ef : errs =          63'b000000000000000000000000000001000000100000000000000000000000000; // D (0x0000000204000000) 
//    12'h37e : errs =          63'b000000000000000000000000000010000000100000000000000000000000000; // D (0x0000000404000000) 
//    12'h85c : errs =          63'b000000000000000000000000000100000000100000000000000000000000000; // D (0x0000000804000000) 
//    12'hb21 : errs =          63'b000000000000000000000000001000000000100000000000000000000000000; // D (0x0000001004000000) 
//    12'hddb : errs =          63'b000000000000000000000000010000000000100000000000000000000000000; // D (0x0000002004000000) 
//    12'h02f : errs =          63'b000000000000000000000000100000000000100000000000000000000000000; // D (0x0000004004000000) 
//    12'hefe : errs =          63'b000000000000000000000001000000000000100000000000000000000000000; // D (0x0000008004000000) 
//    12'h665 : errs =          63'b000000000000000000000010000000000000100000000000000000000000000; // D (0x0000010004000000) 
//    12'h26a : errs =          63'b000000000000000000000100000000000000100000000000000000000000000; // D (0x0000020004000000) 
//    12'ha74 : errs =          63'b000000000000000000001000000000000000100000000000000000000000000; // D (0x0000040004000000) 
//    12'hf71 : errs =          63'b000000000000000000010000000000000000100000000000000000000000000; // D (0x0000080004000000) 
//    12'h57b : errs =          63'b000000000000000000100000000000000000100000000000000000000000000; // D (0x0000100004000000) 
//    12'h456 : errs =          63'b000000000000000001000000000000000000100000000000000000000000000; // D (0x0000200004000000) 
//    12'h60c : errs =          63'b000000000000000010000000000000000000100000000000000000000000000; // D (0x0000400004000000) 
//    12'h2b8 : errs =          63'b000000000000000100000000000000000000100000000000000000000000000; // D (0x0000800004000000) 
//    12'hbd0 : errs =          63'b000000000000001000000000000000000000100000000000000000000000000; // D (0x0001000004000000) 
//    12'hc39 : errs =          63'b000000000000010000000000000000000000100000000000000000000000000; // D (0x0002000004000000) 
//    12'h3eb : errs =          63'b000000000000100000000000000000000000100000000000000000000000000; // D (0x0004000004000000) 
//    12'h976 : errs =          63'b000000000001000000000000000000000000100000000000000000000000000; // D (0x0008000004000000) 
//    12'h975 : errs =          63'b000000000010000000000000000000000000100000000000000000000000000; // D (0x0010000004000000) 
//    12'h973 : errs =          63'b000000000100000000000000000000000000100000000000000000000000000; // D (0x0020000004000000) 
//    12'h97f : errs =          63'b000000001000000000000000000000000000100000000000000000000000000; // D (0x0040000004000000) 
//    12'h967 : errs =          63'b000000010000000000000000000000000000100000000000000000000000000; // D (0x0080000004000000) 
//    12'h957 : errs =          63'b000000100000000000000000000000000000100000000000000000000000000; // D (0x0100000004000000) 
//    12'h937 : errs =          63'b000001000000000000000000000000000000100000000000000000000000000; // D (0x0200000004000000) 
//    12'h9f7 : errs =          63'b000010000000000000000000000000000000100000000000000000000000000; // D (0x0400000004000000) 
//    12'h877 : errs =          63'b000100000000000000000000000000000000100000000000000000000000000; // D (0x0800000004000000) 
//    12'hb77 : errs =          63'b001000000000000000000000000000000000100000000000000000000000000; // D (0x1000000004000000) 
//    12'hd77 : errs =          63'b010000000000000000000000000000000000100000000000000000000000000; // D (0x2000000004000000) 
//    12'h177 : errs =          63'b100000000000000000000000000000000000100000000000000000000000000; // D (0x4000000004000000) 
    12'h2ee : errs =          63'b000000000000000000000000000000000001000000000000000000000000001; // D (0x0000000008000001) 
    12'hda5 : errs =          63'b000000000000000000000000000000000001000000000000000000000000010; // D (0x0000000008000002) 
    12'h60a : errs =          63'b000000000000000000000000000000000001000000000000000000000000100; // D (0x0000000008000004) 
    12'h46d : errs =          63'b000000000000000000000000000000000001000000000000000000000001000; // D (0x0000000008000008) 
    12'h0a3 : errs =          63'b000000000000000000000000000000000001000000000000000000000010000; // D (0x0000000008000010) 
    12'h93f : errs =          63'b000000000000000000000000000000000001000000000000000000000100000; // D (0x0000000008000020) 
    12'hf3e : errs =          63'b000000000000000000000000000000000001000000000000000000001000000; // D (0x0000000008000040) 
    12'h33c : errs =          63'b000000000000000000000000000000000001000000000000000000010000000; // D (0x0000000008000080) 
    12'he01 : errs =          63'b000000000000000000000000000000000001000000000000000000100000000; // D (0x0000000008000100) 
    12'h142 : errs =          63'b000000000000000000000000000000000001000000000000000001000000000; // D (0x0000000008000200) 
    12'hafd : errs =          63'b000000000000000000000000000000000001000000000000000010000000000; // D (0x0000000008000400) 
    12'h8ba : errs =          63'b000000000000000000000000000000000001000000000000000100000000000; // D (0x0000000008000800) 
    12'hc34 : errs =          63'b000000000000000000000000000000000001000000000000001000000000000; // D (0x0000000008001000) 
    12'h528 : errs =          63'b000000000000000000000000000000000001000000000000010000000000000; // D (0x0000000008002000) 
    12'h229 : errs =          63'b000000000000000000000000000000000001000000000000100000000000000; // D (0x0000000008004000) 
    12'hc2b : errs =          63'b000000000000000000000000000000000001000000000001000000000000000; // D (0x0000000008008000) 
    12'h516 : errs =          63'b000000000000000000000000000000000001000000000010000000000000000; // D (0x0000000008010000) 
    12'h255 : errs =          63'b000000000000000000000000000000000001000000000100000000000000000; // D (0x0000000008020000) 
    12'hcd3 : errs =          63'b000000000000000000000000000000000001000000001000000000000000000; // D (0x0000000008040000) 
    12'h4e6 : errs =          63'b000000000000000000000000000000000001000000010000000000000000000; // D (0x0000000008080000) 
    12'h1b5 : errs =          63'b000000000000000000000000000000000001000000100000000000000000000; // D (0x0000000008100000) 
    12'hb13 : errs =          63'b000000000000000000000000000000000001000001000000000000000000000; // D (0x0000000008200000) 
    12'hb66 : errs =          63'b000000000000000000000000000000000001000010000000000000000000000; // D (0x0000000008400000) 
    12'hb8c : errs =          63'b000000000000000000000000000000000001000100000000000000000000000; // D (0x0000000008800000) 
    12'ha58 : errs =          63'b000000000000000000000000000000000001001000000000000000000000000; // D (0x0000000009000000) 
    12'h9f0 : errs =          63'b000000000000000000000000000000000001010000000000000000000000000; // D (0x000000000a000000) 
    12'hea0 : errs =          63'b000000000000000000000000000000000001100000000000000000000000000; // D (0x000000000c000000) 
    12'h7d7 : errs =          63'b000000000000000000000000000000000001000000000000000000000000000; // S (0x0000000008000000) 
//    12'h879 : errs =          63'b000000000000000000000000000000000011000000000000000000000000000; // D (0x0000000018000000) 
//    12'hdb2 : errs =          63'b000000000000000000000000000000000101000000000000000000000000000; // D (0x0000000028000000) 
//    12'h624 : errs =          63'b000000000000000000000000000000001001000000000000000000000000000; // D (0x0000000048000000) 
//    12'h431 : errs =          63'b000000000000000000000000000000010001000000000000000000000000000; // D (0x0000000088000000) 
//    12'h01b : errs =          63'b000000000000000000000000000000100001000000000000000000000000000; // D (0x0000000108000000) 
//    12'h84f : errs =          63'b000000000000000000000000000001000001000000000000000000000000000; // D (0x0000000208000000) 
//    12'hdde : errs =          63'b000000000000000000000000000010000001000000000000000000000000000; // D (0x0000000408000000) 
//    12'h6fc : errs =          63'b000000000000000000000000000100000001000000000000000000000000000; // D (0x0000000808000000) 
//    12'h581 : errs =          63'b000000000000000000000000001000000001000000000000000000000000000; // D (0x0000001008000000) 
//    12'h37b : errs =          63'b000000000000000000000000010000000001000000000000000000000000000; // D (0x0000002008000000) 
//    12'he8f : errs =          63'b000000000000000000000000100000000001000000000000000000000000000; // D (0x0000004008000000) 
//    12'h05e : errs =          63'b000000000000000000000001000000000001000000000000000000000000000; // D (0x0000008008000000) 
//    12'h8c5 : errs =          63'b000000000000000000000010000000000001000000000000000000000000000; // D (0x0000010008000000) 
//    12'hcca : errs =          63'b000000000000000000000100000000000001000000000000000000000000000; // D (0x0000020008000000) 
//    12'h4d4 : errs =          63'b000000000000000000001000000000000001000000000000000000000000000; // D (0x0000040008000000) 
//    12'h1d1 : errs =          63'b000000000000000000010000000000000001000000000000000000000000000; // D (0x0000080008000000) 
//    12'hbdb : errs =          63'b000000000000000000100000000000000001000000000000000000000000000; // D (0x0000100008000000) 
//    12'haf6 : errs =          63'b000000000000000001000000000000000001000000000000000000000000000; // D (0x0000200008000000) 
//    12'h8ac : errs =          63'b000000000000000010000000000000000001000000000000000000000000000; // D (0x0000400008000000) 
//    12'hc18 : errs =          63'b000000000000000100000000000000000001000000000000000000000000000; // D (0x0000800008000000) 
//    12'h570 : errs =          63'b000000000000001000000000000000000001000000000000000000000000000; // D (0x0001000008000000) 
//    12'h299 : errs =          63'b000000000000010000000000000000000001000000000000000000000000000; // D (0x0002000008000000) 
//    12'hd4b : errs =          63'b000000000000100000000000000000000001000000000000000000000000000; // D (0x0004000008000000) 
//    12'h7d6 : errs =          63'b000000000001000000000000000000000001000000000000000000000000000; // D (0x0008000008000000) 
//    12'h7d5 : errs =          63'b000000000010000000000000000000000001000000000000000000000000000; // D (0x0010000008000000) 
//    12'h7d3 : errs =          63'b000000000100000000000000000000000001000000000000000000000000000; // D (0x0020000008000000) 
//    12'h7df : errs =          63'b000000001000000000000000000000000001000000000000000000000000000; // D (0x0040000008000000) 
//    12'h7c7 : errs =          63'b000000010000000000000000000000000001000000000000000000000000000; // D (0x0080000008000000) 
//    12'h7f7 : errs =          63'b000000100000000000000000000000000001000000000000000000000000000; // D (0x0100000008000000) 
//    12'h797 : errs =          63'b000001000000000000000000000000000001000000000000000000000000000; // D (0x0200000008000000) 
//    12'h757 : errs =          63'b000010000000000000000000000000000001000000000000000000000000000; // D (0x0400000008000000) 
//    12'h6d7 : errs =          63'b000100000000000000000000000000000001000000000000000000000000000; // D (0x0800000008000000) 
//    12'h5d7 : errs =          63'b001000000000000000000000000000000001000000000000000000000000000; // D (0x1000000008000000) 
//    12'h3d7 : errs =          63'b010000000000000000000000000000000001000000000000000000000000000; // D (0x2000000008000000) 
//    12'hfd7 : errs =          63'b100000000000000000000000000000000001000000000000000000000000000; // D (0x4000000008000000) 
    12'ha97 : errs =          63'b000000000000000000000000000000000010000000000000000000000000001; // D (0x0000000010000001) 
    12'h5dc : errs =          63'b000000000000000000000000000000000010000000000000000000000000010; // D (0x0000000010000002) 
    12'he73 : errs =          63'b000000000000000000000000000000000010000000000000000000000000100; // D (0x0000000010000004) 
    12'hc14 : errs =          63'b000000000000000000000000000000000010000000000000000000000001000; // D (0x0000000010000008) 
    12'h8da : errs =          63'b000000000000000000000000000000000010000000000000000000000010000; // D (0x0000000010000010) 
    12'h146 : errs =          63'b000000000000000000000000000000000010000000000000000000000100000; // D (0x0000000010000020) 
    12'h747 : errs =          63'b000000000000000000000000000000000010000000000000000000001000000; // D (0x0000000010000040) 
    12'hb45 : errs =          63'b000000000000000000000000000000000010000000000000000000010000000; // D (0x0000000010000080) 
    12'h678 : errs =          63'b000000000000000000000000000000000010000000000000000000100000000; // D (0x0000000010000100) 
    12'h93b : errs =          63'b000000000000000000000000000000000010000000000000000001000000000; // D (0x0000000010000200) 
    12'h284 : errs =          63'b000000000000000000000000000000000010000000000000000010000000000; // D (0x0000000010000400) 
    12'h0c3 : errs =          63'b000000000000000000000000000000000010000000000000000100000000000; // D (0x0000000010000800) 
    12'h44d : errs =          63'b000000000000000000000000000000000010000000000000001000000000000; // D (0x0000000010001000) 
    12'hd51 : errs =          63'b000000000000000000000000000000000010000000000000010000000000000; // D (0x0000000010002000) 
    12'ha50 : errs =          63'b000000000000000000000000000000000010000000000000100000000000000; // D (0x0000000010004000) 
    12'h452 : errs =          63'b000000000000000000000000000000000010000000000001000000000000000; // D (0x0000000010008000) 
    12'hd6f : errs =          63'b000000000000000000000000000000000010000000000010000000000000000; // D (0x0000000010010000) 
    12'ha2c : errs =          63'b000000000000000000000000000000000010000000000100000000000000000; // D (0x0000000010020000) 
    12'h4aa : errs =          63'b000000000000000000000000000000000010000000001000000000000000000; // D (0x0000000010040000) 
    12'hc9f : errs =          63'b000000000000000000000000000000000010000000010000000000000000000; // D (0x0000000010080000) 
    12'h9cc : errs =          63'b000000000000000000000000000000000010000000100000000000000000000; // D (0x0000000010100000) 
    12'h36a : errs =          63'b000000000000000000000000000000000010000001000000000000000000000; // D (0x0000000010200000) 
    12'h31f : errs =          63'b000000000000000000000000000000000010000010000000000000000000000; // D (0x0000000010400000) 
    12'h3f5 : errs =          63'b000000000000000000000000000000000010000100000000000000000000000; // D (0x0000000010800000) 
    12'h221 : errs =          63'b000000000000000000000000000000000010001000000000000000000000000; // D (0x0000000011000000) 
    12'h189 : errs =          63'b000000000000000000000000000000000010010000000000000000000000000; // D (0x0000000012000000) 
    12'h6d9 : errs =          63'b000000000000000000000000000000000010100000000000000000000000000; // D (0x0000000014000000) 
    12'h879 : errs =          63'b000000000000000000000000000000000011000000000000000000000000000; // D (0x0000000018000000) 
    12'hfae : errs =          63'b000000000000000000000000000000000010000000000000000000000000000; // S (0x0000000010000000) 
//    12'h5cb : errs =          63'b000000000000000000000000000000000110000000000000000000000000000; // D (0x0000000030000000) 
//    12'he5d : errs =          63'b000000000000000000000000000000001010000000000000000000000000000; // D (0x0000000050000000) 
//    12'hc48 : errs =          63'b000000000000000000000000000000010010000000000000000000000000000; // D (0x0000000090000000) 
//    12'h862 : errs =          63'b000000000000000000000000000000100010000000000000000000000000000; // D (0x0000000110000000) 
//    12'h036 : errs =          63'b000000000000000000000000000001000010000000000000000000000000000; // D (0x0000000210000000) 
//    12'h5a7 : errs =          63'b000000000000000000000000000010000010000000000000000000000000000; // D (0x0000000410000000) 
//    12'he85 : errs =          63'b000000000000000000000000000100000010000000000000000000000000000; // D (0x0000000810000000) 
//    12'hdf8 : errs =          63'b000000000000000000000000001000000010000000000000000000000000000; // D (0x0000001010000000) 
//    12'hb02 : errs =          63'b000000000000000000000000010000000010000000000000000000000000000; // D (0x0000002010000000) 
//    12'h6f6 : errs =          63'b000000000000000000000000100000000010000000000000000000000000000; // D (0x0000004010000000) 
//    12'h827 : errs =          63'b000000000000000000000001000000000010000000000000000000000000000; // D (0x0000008010000000) 
//    12'h0bc : errs =          63'b000000000000000000000010000000000010000000000000000000000000000; // D (0x0000010010000000) 
//    12'h4b3 : errs =          63'b000000000000000000000100000000000010000000000000000000000000000; // D (0x0000020010000000) 
//    12'hcad : errs =          63'b000000000000000000001000000000000010000000000000000000000000000; // D (0x0000040010000000) 
//    12'h9a8 : errs =          63'b000000000000000000010000000000000010000000000000000000000000000; // D (0x0000080010000000) 
//    12'h3a2 : errs =          63'b000000000000000000100000000000000010000000000000000000000000000; // D (0x0000100010000000) 
//    12'h28f : errs =          63'b000000000000000001000000000000000010000000000000000000000000000; // D (0x0000200010000000) 
//    12'h0d5 : errs =          63'b000000000000000010000000000000000010000000000000000000000000000; // D (0x0000400010000000) 
//    12'h461 : errs =          63'b000000000000000100000000000000000010000000000000000000000000000; // D (0x0000800010000000) 
//    12'hd09 : errs =          63'b000000000000001000000000000000000010000000000000000000000000000; // D (0x0001000010000000) 
//    12'hae0 : errs =          63'b000000000000010000000000000000000010000000000000000000000000000; // D (0x0002000010000000) 
//    12'h532 : errs =          63'b000000000000100000000000000000000010000000000000000000000000000; // D (0x0004000010000000) 
//    12'hfaf : errs =          63'b000000000001000000000000000000000010000000000000000000000000000; // D (0x0008000010000000) 
//    12'hfac : errs =          63'b000000000010000000000000000000000010000000000000000000000000000; // D (0x0010000010000000) 
//    12'hfaa : errs =          63'b000000000100000000000000000000000010000000000000000000000000000; // D (0x0020000010000000) 
//    12'hfa6 : errs =          63'b000000001000000000000000000000000010000000000000000000000000000; // D (0x0040000010000000) 
//    12'hfbe : errs =          63'b000000010000000000000000000000000010000000000000000000000000000; // D (0x0080000010000000) 
//    12'hf8e : errs =          63'b000000100000000000000000000000000010000000000000000000000000000; // D (0x0100000010000000) 
//    12'hfee : errs =          63'b000001000000000000000000000000000010000000000000000000000000000; // D (0x0200000010000000) 
//    12'hf2e : errs =          63'b000010000000000000000000000000000010000000000000000000000000000; // D (0x0400000010000000) 
//    12'heae : errs =          63'b000100000000000000000000000000000010000000000000000000000000000; // D (0x0800000010000000) 
//    12'hdae : errs =          63'b001000000000000000000000000000000010000000000000000000000000000; // D (0x1000000010000000) 
//    12'hbae : errs =          63'b010000000000000000000000000000000010000000000000000000000000000; // D (0x2000000010000000) 
//    12'h7ae : errs =          63'b100000000000000000000000000000000010000000000000000000000000000; // D (0x4000000010000000) 
    12'hf5c : errs =          63'b000000000000000000000000000000000100000000000000000000000000001; // D (0x0000000020000001) 
    12'h017 : errs =          63'b000000000000000000000000000000000100000000000000000000000000010; // D (0x0000000020000002) 
    12'hbb8 : errs =          63'b000000000000000000000000000000000100000000000000000000000000100; // D (0x0000000020000004) 
    12'h9df : errs =          63'b000000000000000000000000000000000100000000000000000000000001000; // D (0x0000000020000008) 
    12'hd11 : errs =          63'b000000000000000000000000000000000100000000000000000000000010000; // D (0x0000000020000010) 
    12'h48d : errs =          63'b000000000000000000000000000000000100000000000000000000000100000; // D (0x0000000020000020) 
    12'h28c : errs =          63'b000000000000000000000000000000000100000000000000000000001000000; // D (0x0000000020000040) 
    12'he8e : errs =          63'b000000000000000000000000000000000100000000000000000000010000000; // D (0x0000000020000080) 
    12'h3b3 : errs =          63'b000000000000000000000000000000000100000000000000000000100000000; // D (0x0000000020000100) 
    12'hcf0 : errs =          63'b000000000000000000000000000000000100000000000000000001000000000; // D (0x0000000020000200) 
    12'h74f : errs =          63'b000000000000000000000000000000000100000000000000000010000000000; // D (0x0000000020000400) 
    12'h508 : errs =          63'b000000000000000000000000000000000100000000000000000100000000000; // D (0x0000000020000800) 
    12'h186 : errs =          63'b000000000000000000000000000000000100000000000000001000000000000; // D (0x0000000020001000) 
    12'h89a : errs =          63'b000000000000000000000000000000000100000000000000010000000000000; // D (0x0000000020002000) 
    12'hf9b : errs =          63'b000000000000000000000000000000000100000000000000100000000000000; // D (0x0000000020004000) 
    12'h199 : errs =          63'b000000000000000000000000000000000100000000000001000000000000000; // D (0x0000000020008000) 
    12'h8a4 : errs =          63'b000000000000000000000000000000000100000000000010000000000000000; // D (0x0000000020010000) 
    12'hfe7 : errs =          63'b000000000000000000000000000000000100000000000100000000000000000; // D (0x0000000020020000) 
    12'h161 : errs =          63'b000000000000000000000000000000000100000000001000000000000000000; // D (0x0000000020040000) 
    12'h954 : errs =          63'b000000000000000000000000000000000100000000010000000000000000000; // D (0x0000000020080000) 
    12'hc07 : errs =          63'b000000000000000000000000000000000100000000100000000000000000000; // D (0x0000000020100000) 
    12'h6a1 : errs =          63'b000000000000000000000000000000000100000001000000000000000000000; // D (0x0000000020200000) 
    12'h6d4 : errs =          63'b000000000000000000000000000000000100000010000000000000000000000; // D (0x0000000020400000) 
    12'h63e : errs =          63'b000000000000000000000000000000000100000100000000000000000000000; // D (0x0000000020800000) 
    12'h7ea : errs =          63'b000000000000000000000000000000000100001000000000000000000000000; // D (0x0000000021000000) 
    12'h442 : errs =          63'b000000000000000000000000000000000100010000000000000000000000000; // D (0x0000000022000000) 
    12'h312 : errs =          63'b000000000000000000000000000000000100100000000000000000000000000; // D (0x0000000024000000) 
    12'hdb2 : errs =          63'b000000000000000000000000000000000101000000000000000000000000000; // D (0x0000000028000000) 
    12'h5cb : errs =          63'b000000000000000000000000000000000110000000000000000000000000000; // D (0x0000000030000000) 
    12'ha65 : errs =          63'b000000000000000000000000000000000100000000000000000000000000000; // S (0x0000000020000000) 
//    12'hb96 : errs =          63'b000000000000000000000000000000001100000000000000000000000000000; // D (0x0000000060000000) 
//    12'h983 : errs =          63'b000000000000000000000000000000010100000000000000000000000000000; // D (0x00000000a0000000) 
//    12'hda9 : errs =          63'b000000000000000000000000000000100100000000000000000000000000000; // D (0x0000000120000000) 
//    12'h5fd : errs =          63'b000000000000000000000000000001000100000000000000000000000000000; // D (0x0000000220000000) 
//    12'h06c : errs =          63'b000000000000000000000000000010000100000000000000000000000000000; // D (0x0000000420000000) 
//    12'hb4e : errs =          63'b000000000000000000000000000100000100000000000000000000000000000; // D (0x0000000820000000) 
//    12'h833 : errs =          63'b000000000000000000000000001000000100000000000000000000000000000; // D (0x0000001020000000) 
//    12'hec9 : errs =          63'b000000000000000000000000010000000100000000000000000000000000000; // D (0x0000002020000000) 
//    12'h33d : errs =          63'b000000000000000000000000100000000100000000000000000000000000000; // D (0x0000004020000000) 
//    12'hdec : errs =          63'b000000000000000000000001000000000100000000000000000000000000000; // D (0x0000008020000000) 
//    12'h577 : errs =          63'b000000000000000000000010000000000100000000000000000000000000000; // D (0x0000010020000000) 
//    12'h178 : errs =          63'b000000000000000000000100000000000100000000000000000000000000000; // D (0x0000020020000000) 
//    12'h966 : errs =          63'b000000000000000000001000000000000100000000000000000000000000000; // D (0x0000040020000000) 
//    12'hc63 : errs =          63'b000000000000000000010000000000000100000000000000000000000000000; // D (0x0000080020000000) 
//    12'h669 : errs =          63'b000000000000000000100000000000000100000000000000000000000000000; // D (0x0000100020000000) 
//    12'h744 : errs =          63'b000000000000000001000000000000000100000000000000000000000000000; // D (0x0000200020000000) 
//    12'h51e : errs =          63'b000000000000000010000000000000000100000000000000000000000000000; // D (0x0000400020000000) 
//    12'h1aa : errs =          63'b000000000000000100000000000000000100000000000000000000000000000; // D (0x0000800020000000) 
//    12'h8c2 : errs =          63'b000000000000001000000000000000000100000000000000000000000000000; // D (0x0001000020000000) 
//    12'hf2b : errs =          63'b000000000000010000000000000000000100000000000000000000000000000; // D (0x0002000020000000) 
//    12'h0f9 : errs =          63'b000000000000100000000000000000000100000000000000000000000000000; // D (0x0004000020000000) 
//    12'ha64 : errs =          63'b000000000001000000000000000000000100000000000000000000000000000; // D (0x0008000020000000) 
//    12'ha67 : errs =          63'b000000000010000000000000000000000100000000000000000000000000000; // D (0x0010000020000000) 
//    12'ha61 : errs =          63'b000000000100000000000000000000000100000000000000000000000000000; // D (0x0020000020000000) 
//    12'ha6d : errs =          63'b000000001000000000000000000000000100000000000000000000000000000; // D (0x0040000020000000) 
//    12'ha75 : errs =          63'b000000010000000000000000000000000100000000000000000000000000000; // D (0x0080000020000000) 
//    12'ha45 : errs =          63'b000000100000000000000000000000000100000000000000000000000000000; // D (0x0100000020000000) 
//    12'ha25 : errs =          63'b000001000000000000000000000000000100000000000000000000000000000; // D (0x0200000020000000) 
//    12'hae5 : errs =          63'b000010000000000000000000000000000100000000000000000000000000000; // D (0x0400000020000000) 
//    12'hb65 : errs =          63'b000100000000000000000000000000000100000000000000000000000000000; // D (0x0800000020000000) 
//    12'h865 : errs =          63'b001000000000000000000000000000000100000000000000000000000000000; // D (0x1000000020000000) 
//    12'he65 : errs =          63'b010000000000000000000000000000000100000000000000000000000000000; // D (0x2000000020000000) 
//    12'h265 : errs =          63'b100000000000000000000000000000000100000000000000000000000000000; // D (0x4000000020000000) 
    12'h4ca : errs =          63'b000000000000000000000000000000001000000000000000000000000000001; // D (0x0000000040000001) 
    12'hb81 : errs =          63'b000000000000000000000000000000001000000000000000000000000000010; // D (0x0000000040000002) 
    12'h02e : errs =          63'b000000000000000000000000000000001000000000000000000000000000100; // D (0x0000000040000004) 
    12'h249 : errs =          63'b000000000000000000000000000000001000000000000000000000000001000; // D (0x0000000040000008) 
    12'h687 : errs =          63'b000000000000000000000000000000001000000000000000000000000010000; // D (0x0000000040000010) 
    12'hf1b : errs =          63'b000000000000000000000000000000001000000000000000000000000100000; // D (0x0000000040000020) 
    12'h91a : errs =          63'b000000000000000000000000000000001000000000000000000000001000000; // D (0x0000000040000040) 
    12'h518 : errs =          63'b000000000000000000000000000000001000000000000000000000010000000; // D (0x0000000040000080) 
    12'h825 : errs =          63'b000000000000000000000000000000001000000000000000000000100000000; // D (0x0000000040000100) 
    12'h766 : errs =          63'b000000000000000000000000000000001000000000000000000001000000000; // D (0x0000000040000200) 
    12'hcd9 : errs =          63'b000000000000000000000000000000001000000000000000000010000000000; // D (0x0000000040000400) 
    12'he9e : errs =          63'b000000000000000000000000000000001000000000000000000100000000000; // D (0x0000000040000800) 
    12'ha10 : errs =          63'b000000000000000000000000000000001000000000000000001000000000000; // D (0x0000000040001000) 
    12'h30c : errs =          63'b000000000000000000000000000000001000000000000000010000000000000; // D (0x0000000040002000) 
    12'h40d : errs =          63'b000000000000000000000000000000001000000000000000100000000000000; // D (0x0000000040004000) 
    12'ha0f : errs =          63'b000000000000000000000000000000001000000000000001000000000000000; // D (0x0000000040008000) 
    12'h332 : errs =          63'b000000000000000000000000000000001000000000000010000000000000000; // D (0x0000000040010000) 
    12'h471 : errs =          63'b000000000000000000000000000000001000000000000100000000000000000; // D (0x0000000040020000) 
    12'haf7 : errs =          63'b000000000000000000000000000000001000000000001000000000000000000; // D (0x0000000040040000) 
    12'h2c2 : errs =          63'b000000000000000000000000000000001000000000010000000000000000000; // D (0x0000000040080000) 
    12'h791 : errs =          63'b000000000000000000000000000000001000000000100000000000000000000; // D (0x0000000040100000) 
    12'hd37 : errs =          63'b000000000000000000000000000000001000000001000000000000000000000; // D (0x0000000040200000) 
    12'hd42 : errs =          63'b000000000000000000000000000000001000000010000000000000000000000; // D (0x0000000040400000) 
    12'hda8 : errs =          63'b000000000000000000000000000000001000000100000000000000000000000; // D (0x0000000040800000) 
    12'hc7c : errs =          63'b000000000000000000000000000000001000001000000000000000000000000; // D (0x0000000041000000) 
    12'hfd4 : errs =          63'b000000000000000000000000000000001000010000000000000000000000000; // D (0x0000000042000000) 
    12'h884 : errs =          63'b000000000000000000000000000000001000100000000000000000000000000; // D (0x0000000044000000) 
    12'h624 : errs =          63'b000000000000000000000000000000001001000000000000000000000000000; // D (0x0000000048000000) 
    12'he5d : errs =          63'b000000000000000000000000000000001010000000000000000000000000000; // D (0x0000000050000000) 
    12'hb96 : errs =          63'b000000000000000000000000000000001100000000000000000000000000000; // D (0x0000000060000000) 
    12'h1f3 : errs =          63'b000000000000000000000000000000001000000000000000000000000000000; // S (0x0000000040000000) 
//    12'h215 : errs =          63'b000000000000000000000000000000011000000000000000000000000000000; // D (0x00000000c0000000) 
//    12'h63f : errs =          63'b000000000000000000000000000000101000000000000000000000000000000; // D (0x0000000140000000) 
//    12'he6b : errs =          63'b000000000000000000000000000001001000000000000000000000000000000; // D (0x0000000240000000) 
//    12'hbfa : errs =          63'b000000000000000000000000000010001000000000000000000000000000000; // D (0x0000000440000000) 
//    12'h0d8 : errs =          63'b000000000000000000000000000100001000000000000000000000000000000; // D (0x0000000840000000) 
//    12'h3a5 : errs =          63'b000000000000000000000000001000001000000000000000000000000000000; // D (0x0000001040000000) 
//    12'h55f : errs =          63'b000000000000000000000000010000001000000000000000000000000000000; // D (0x0000002040000000) 
//    12'h8ab : errs =          63'b000000000000000000000000100000001000000000000000000000000000000; // D (0x0000004040000000) 
//    12'h67a : errs =          63'b000000000000000000000001000000001000000000000000000000000000000; // D (0x0000008040000000) 
//    12'hee1 : errs =          63'b000000000000000000000010000000001000000000000000000000000000000; // D (0x0000010040000000) 
//    12'haee : errs =          63'b000000000000000000000100000000001000000000000000000000000000000; // D (0x0000020040000000) 
//    12'h2f0 : errs =          63'b000000000000000000001000000000001000000000000000000000000000000; // D (0x0000040040000000) 
//    12'h7f5 : errs =          63'b000000000000000000010000000000001000000000000000000000000000000; // D (0x0000080040000000) 
//    12'hdff : errs =          63'b000000000000000000100000000000001000000000000000000000000000000; // D (0x0000100040000000) 
//    12'hcd2 : errs =          63'b000000000000000001000000000000001000000000000000000000000000000; // D (0x0000200040000000) 
//    12'he88 : errs =          63'b000000000000000010000000000000001000000000000000000000000000000; // D (0x0000400040000000) 
//    12'ha3c : errs =          63'b000000000000000100000000000000001000000000000000000000000000000; // D (0x0000800040000000) 
//    12'h354 : errs =          63'b000000000000001000000000000000001000000000000000000000000000000; // D (0x0001000040000000) 
//    12'h4bd : errs =          63'b000000000000010000000000000000001000000000000000000000000000000; // D (0x0002000040000000) 
//    12'hb6f : errs =          63'b000000000000100000000000000000001000000000000000000000000000000; // D (0x0004000040000000) 
//    12'h1f2 : errs =          63'b000000000001000000000000000000001000000000000000000000000000000; // D (0x0008000040000000) 
//    12'h1f1 : errs =          63'b000000000010000000000000000000001000000000000000000000000000000; // D (0x0010000040000000) 
//    12'h1f7 : errs =          63'b000000000100000000000000000000001000000000000000000000000000000; // D (0x0020000040000000) 
//    12'h1fb : errs =          63'b000000001000000000000000000000001000000000000000000000000000000; // D (0x0040000040000000) 
//    12'h1e3 : errs =          63'b000000010000000000000000000000001000000000000000000000000000000; // D (0x0080000040000000) 
//    12'h1d3 : errs =          63'b000000100000000000000000000000001000000000000000000000000000000; // D (0x0100000040000000) 
//    12'h1b3 : errs =          63'b000001000000000000000000000000001000000000000000000000000000000; // D (0x0200000040000000) 
//    12'h173 : errs =          63'b000010000000000000000000000000001000000000000000000000000000000; // D (0x0400000040000000) 
//    12'h0f3 : errs =          63'b000100000000000000000000000000001000000000000000000000000000000; // D (0x0800000040000000) 
//    12'h3f3 : errs =          63'b001000000000000000000000000000001000000000000000000000000000000; // D (0x1000000040000000) 
//    12'h5f3 : errs =          63'b010000000000000000000000000000001000000000000000000000000000000; // D (0x2000000040000000) 
//    12'h9f3 : errs =          63'b100000000000000000000000000000001000000000000000000000000000000; // D (0x4000000040000000) 
    12'h6df : errs =          63'b000000000000000000000000000000010000000000000000000000000000001; // D (0x0000000080000001) 
    12'h994 : errs =          63'b000000000000000000000000000000010000000000000000000000000000010; // D (0x0000000080000002) 
    12'h23b : errs =          63'b000000000000000000000000000000010000000000000000000000000000100; // D (0x0000000080000004) 
    12'h05c : errs =          63'b000000000000000000000000000000010000000000000000000000000001000; // D (0x0000000080000008) 
    12'h492 : errs =          63'b000000000000000000000000000000010000000000000000000000000010000; // D (0x0000000080000010) 
    12'hd0e : errs =          63'b000000000000000000000000000000010000000000000000000000000100000; // D (0x0000000080000020) 
    12'hb0f : errs =          63'b000000000000000000000000000000010000000000000000000000001000000; // D (0x0000000080000040) 
    12'h70d : errs =          63'b000000000000000000000000000000010000000000000000000000010000000; // D (0x0000000080000080) 
    12'ha30 : errs =          63'b000000000000000000000000000000010000000000000000000000100000000; // D (0x0000000080000100) 
    12'h573 : errs =          63'b000000000000000000000000000000010000000000000000000001000000000; // D (0x0000000080000200) 
    12'hecc : errs =          63'b000000000000000000000000000000010000000000000000000010000000000; // D (0x0000000080000400) 
    12'hc8b : errs =          63'b000000000000000000000000000000010000000000000000000100000000000; // D (0x0000000080000800) 
    12'h805 : errs =          63'b000000000000000000000000000000010000000000000000001000000000000; // D (0x0000000080001000) 
    12'h119 : errs =          63'b000000000000000000000000000000010000000000000000010000000000000; // D (0x0000000080002000) 
    12'h618 : errs =          63'b000000000000000000000000000000010000000000000000100000000000000; // D (0x0000000080004000) 
    12'h81a : errs =          63'b000000000000000000000000000000010000000000000001000000000000000; // D (0x0000000080008000) 
    12'h127 : errs =          63'b000000000000000000000000000000010000000000000010000000000000000; // D (0x0000000080010000) 
    12'h664 : errs =          63'b000000000000000000000000000000010000000000000100000000000000000; // D (0x0000000080020000) 
    12'h8e2 : errs =          63'b000000000000000000000000000000010000000000001000000000000000000; // D (0x0000000080040000) 
    12'h0d7 : errs =          63'b000000000000000000000000000000010000000000010000000000000000000; // D (0x0000000080080000) 
    12'h584 : errs =          63'b000000000000000000000000000000010000000000100000000000000000000; // D (0x0000000080100000) 
    12'hf22 : errs =          63'b000000000000000000000000000000010000000001000000000000000000000; // D (0x0000000080200000) 
    12'hf57 : errs =          63'b000000000000000000000000000000010000000010000000000000000000000; // D (0x0000000080400000) 
    12'hfbd : errs =          63'b000000000000000000000000000000010000000100000000000000000000000; // D (0x0000000080800000) 
    12'he69 : errs =          63'b000000000000000000000000000000010000001000000000000000000000000; // D (0x0000000081000000) 
    12'hdc1 : errs =          63'b000000000000000000000000000000010000010000000000000000000000000; // D (0x0000000082000000) 
    12'ha91 : errs =          63'b000000000000000000000000000000010000100000000000000000000000000; // D (0x0000000084000000) 
    12'h431 : errs =          63'b000000000000000000000000000000010001000000000000000000000000000; // D (0x0000000088000000) 
    12'hc48 : errs =          63'b000000000000000000000000000000010010000000000000000000000000000; // D (0x0000000090000000) 
    12'h983 : errs =          63'b000000000000000000000000000000010100000000000000000000000000000; // D (0x00000000a0000000) 
    12'h215 : errs =          63'b000000000000000000000000000000011000000000000000000000000000000; // D (0x00000000c0000000) 
    12'h3e6 : errs =          63'b000000000000000000000000000000010000000000000000000000000000000; // S (0x0000000080000000) 
//    12'h42a : errs =          63'b000000000000000000000000000000110000000000000000000000000000000; // D (0x0000000180000000) 
//    12'hc7e : errs =          63'b000000000000000000000000000001010000000000000000000000000000000; // D (0x0000000280000000) 
//    12'h9ef : errs =          63'b000000000000000000000000000010010000000000000000000000000000000; // D (0x0000000480000000) 
//    12'h2cd : errs =          63'b000000000000000000000000000100010000000000000000000000000000000; // D (0x0000000880000000) 
//    12'h1b0 : errs =          63'b000000000000000000000000001000010000000000000000000000000000000; // D (0x0000001080000000) 
//    12'h74a : errs =          63'b000000000000000000000000010000010000000000000000000000000000000; // D (0x0000002080000000) 
//    12'habe : errs =          63'b000000000000000000000000100000010000000000000000000000000000000; // D (0x0000004080000000) 
//    12'h46f : errs =          63'b000000000000000000000001000000010000000000000000000000000000000; // D (0x0000008080000000) 
//    12'hcf4 : errs =          63'b000000000000000000000010000000010000000000000000000000000000000; // D (0x0000010080000000) 
//    12'h8fb : errs =          63'b000000000000000000000100000000010000000000000000000000000000000; // D (0x0000020080000000) 
//    12'h0e5 : errs =          63'b000000000000000000001000000000010000000000000000000000000000000; // D (0x0000040080000000) 
//    12'h5e0 : errs =          63'b000000000000000000010000000000010000000000000000000000000000000; // D (0x0000080080000000) 
//    12'hfea : errs =          63'b000000000000000000100000000000010000000000000000000000000000000; // D (0x0000100080000000) 
//    12'hec7 : errs =          63'b000000000000000001000000000000010000000000000000000000000000000; // D (0x0000200080000000) 
//    12'hc9d : errs =          63'b000000000000000010000000000000010000000000000000000000000000000; // D (0x0000400080000000) 
//    12'h829 : errs =          63'b000000000000000100000000000000010000000000000000000000000000000; // D (0x0000800080000000) 
//    12'h141 : errs =          63'b000000000000001000000000000000010000000000000000000000000000000; // D (0x0001000080000000) 
//    12'h6a8 : errs =          63'b000000000000010000000000000000010000000000000000000000000000000; // D (0x0002000080000000) 
//    12'h97a : errs =          63'b000000000000100000000000000000010000000000000000000000000000000; // D (0x0004000080000000) 
//    12'h3e7 : errs =          63'b000000000001000000000000000000010000000000000000000000000000000; // D (0x0008000080000000) 
//    12'h3e4 : errs =          63'b000000000010000000000000000000010000000000000000000000000000000; // D (0x0010000080000000) 
//    12'h3e2 : errs =          63'b000000000100000000000000000000010000000000000000000000000000000; // D (0x0020000080000000) 
//    12'h3ee : errs =          63'b000000001000000000000000000000010000000000000000000000000000000; // D (0x0040000080000000) 
//    12'h3f6 : errs =          63'b000000010000000000000000000000010000000000000000000000000000000; // D (0x0080000080000000) 
//    12'h3c6 : errs =          63'b000000100000000000000000000000010000000000000000000000000000000; // D (0x0100000080000000) 
//    12'h3a6 : errs =          63'b000001000000000000000000000000010000000000000000000000000000000; // D (0x0200000080000000) 
//    12'h366 : errs =          63'b000010000000000000000000000000010000000000000000000000000000000; // D (0x0400000080000000) 
//    12'h2e6 : errs =          63'b000100000000000000000000000000010000000000000000000000000000000; // D (0x0800000080000000) 
//    12'h1e6 : errs =          63'b001000000000000000000000000000010000000000000000000000000000000; // D (0x1000000080000000) 
//    12'h7e6 : errs =          63'b010000000000000000000000000000010000000000000000000000000000000; // D (0x2000000080000000) 
//    12'hbe6 : errs =          63'b100000000000000000000000000000010000000000000000000000000000000; // D (0x4000000080000000) 
    12'h2f5 : errs =          63'b000000000000000000000000000000100000000000000000000000000000001; // D (0x0000000100000001) 
    12'hdbe : errs =          63'b000000000000000000000000000000100000000000000000000000000000010; // D (0x0000000100000002) 
    12'h611 : errs =          63'b000000000000000000000000000000100000000000000000000000000000100; // D (0x0000000100000004) 
    12'h476 : errs =          63'b000000000000000000000000000000100000000000000000000000000001000; // D (0x0000000100000008) 
    12'h0b8 : errs =          63'b000000000000000000000000000000100000000000000000000000000010000; // D (0x0000000100000010) 
    12'h924 : errs =          63'b000000000000000000000000000000100000000000000000000000000100000; // D (0x0000000100000020) 
    12'hf25 : errs =          63'b000000000000000000000000000000100000000000000000000000001000000; // D (0x0000000100000040) 
    12'h327 : errs =          63'b000000000000000000000000000000100000000000000000000000010000000; // D (0x0000000100000080) 
    12'he1a : errs =          63'b000000000000000000000000000000100000000000000000000000100000000; // D (0x0000000100000100) 
    12'h159 : errs =          63'b000000000000000000000000000000100000000000000000000001000000000; // D (0x0000000100000200) 
    12'hae6 : errs =          63'b000000000000000000000000000000100000000000000000000010000000000; // D (0x0000000100000400) 
    12'h8a1 : errs =          63'b000000000000000000000000000000100000000000000000000100000000000; // D (0x0000000100000800) 
    12'hc2f : errs =          63'b000000000000000000000000000000100000000000000000001000000000000; // D (0x0000000100001000) 
    12'h533 : errs =          63'b000000000000000000000000000000100000000000000000010000000000000; // D (0x0000000100002000) 
    12'h232 : errs =          63'b000000000000000000000000000000100000000000000000100000000000000; // D (0x0000000100004000) 
    12'hc30 : errs =          63'b000000000000000000000000000000100000000000000001000000000000000; // D (0x0000000100008000) 
    12'h50d : errs =          63'b000000000000000000000000000000100000000000000010000000000000000; // D (0x0000000100010000) 
    12'h24e : errs =          63'b000000000000000000000000000000100000000000000100000000000000000; // D (0x0000000100020000) 
    12'hcc8 : errs =          63'b000000000000000000000000000000100000000000001000000000000000000; // D (0x0000000100040000) 
    12'h4fd : errs =          63'b000000000000000000000000000000100000000000010000000000000000000; // D (0x0000000100080000) 
    12'h1ae : errs =          63'b000000000000000000000000000000100000000000100000000000000000000; // D (0x0000000100100000) 
    12'hb08 : errs =          63'b000000000000000000000000000000100000000001000000000000000000000; // D (0x0000000100200000) 
    12'hb7d : errs =          63'b000000000000000000000000000000100000000010000000000000000000000; // D (0x0000000100400000) 
    12'hb97 : errs =          63'b000000000000000000000000000000100000000100000000000000000000000; // D (0x0000000100800000) 
    12'ha43 : errs =          63'b000000000000000000000000000000100000001000000000000000000000000; // D (0x0000000101000000) 
    12'h9eb : errs =          63'b000000000000000000000000000000100000010000000000000000000000000; // D (0x0000000102000000) 
    12'hebb : errs =          63'b000000000000000000000000000000100000100000000000000000000000000; // D (0x0000000104000000) 
    12'h01b : errs =          63'b000000000000000000000000000000100001000000000000000000000000000; // D (0x0000000108000000) 
    12'h862 : errs =          63'b000000000000000000000000000000100010000000000000000000000000000; // D (0x0000000110000000) 
    12'hda9 : errs =          63'b000000000000000000000000000000100100000000000000000000000000000; // D (0x0000000120000000) 
    12'h63f : errs =          63'b000000000000000000000000000000101000000000000000000000000000000; // D (0x0000000140000000) 
    12'h42a : errs =          63'b000000000000000000000000000000110000000000000000000000000000000; // D (0x0000000180000000) 
    12'h7cc : errs =          63'b000000000000000000000000000000100000000000000000000000000000000; // S (0x0000000100000000) 
//    12'h854 : errs =          63'b000000000000000000000000000001100000000000000000000000000000000; // D (0x0000000300000000) 
//    12'hdc5 : errs =          63'b000000000000000000000000000010100000000000000000000000000000000; // D (0x0000000500000000) 
//    12'h6e7 : errs =          63'b000000000000000000000000000100100000000000000000000000000000000; // D (0x0000000900000000) 
//    12'h59a : errs =          63'b000000000000000000000000001000100000000000000000000000000000000; // D (0x0000001100000000) 
//    12'h360 : errs =          63'b000000000000000000000000010000100000000000000000000000000000000; // D (0x0000002100000000) 
//    12'he94 : errs =          63'b000000000000000000000000100000100000000000000000000000000000000; // D (0x0000004100000000) 
//    12'h045 : errs =          63'b000000000000000000000001000000100000000000000000000000000000000; // D (0x0000008100000000) 
//    12'h8de : errs =          63'b000000000000000000000010000000100000000000000000000000000000000; // D (0x0000010100000000) 
//    12'hcd1 : errs =          63'b000000000000000000000100000000100000000000000000000000000000000; // D (0x0000020100000000) 
//    12'h4cf : errs =          63'b000000000000000000001000000000100000000000000000000000000000000; // D (0x0000040100000000) 
//    12'h1ca : errs =          63'b000000000000000000010000000000100000000000000000000000000000000; // D (0x0000080100000000) 
//    12'hbc0 : errs =          63'b000000000000000000100000000000100000000000000000000000000000000; // D (0x0000100100000000) 
//    12'haed : errs =          63'b000000000000000001000000000000100000000000000000000000000000000; // D (0x0000200100000000) 
//    12'h8b7 : errs =          63'b000000000000000010000000000000100000000000000000000000000000000; // D (0x0000400100000000) 
//    12'hc03 : errs =          63'b000000000000000100000000000000100000000000000000000000000000000; // D (0x0000800100000000) 
//    12'h56b : errs =          63'b000000000000001000000000000000100000000000000000000000000000000; // D (0x0001000100000000) 
//    12'h282 : errs =          63'b000000000000010000000000000000100000000000000000000000000000000; // D (0x0002000100000000) 
//    12'hd50 : errs =          63'b000000000000100000000000000000100000000000000000000000000000000; // D (0x0004000100000000) 
//    12'h7cd : errs =          63'b000000000001000000000000000000100000000000000000000000000000000; // D (0x0008000100000000) 
//    12'h7ce : errs =          63'b000000000010000000000000000000100000000000000000000000000000000; // D (0x0010000100000000) 
//    12'h7c8 : errs =          63'b000000000100000000000000000000100000000000000000000000000000000; // D (0x0020000100000000) 
//    12'h7c4 : errs =          63'b000000001000000000000000000000100000000000000000000000000000000; // D (0x0040000100000000) 
//    12'h7dc : errs =          63'b000000010000000000000000000000100000000000000000000000000000000; // D (0x0080000100000000) 
//    12'h7ec : errs =          63'b000000100000000000000000000000100000000000000000000000000000000; // D (0x0100000100000000) 
//    12'h78c : errs =          63'b000001000000000000000000000000100000000000000000000000000000000; // D (0x0200000100000000) 
//    12'h74c : errs =          63'b000010000000000000000000000000100000000000000000000000000000000; // D (0x0400000100000000) 
//    12'h6cc : errs =          63'b000100000000000000000000000000100000000000000000000000000000000; // D (0x0800000100000000) 
//    12'h5cc : errs =          63'b001000000000000000000000000000100000000000000000000000000000000; // D (0x1000000100000000) 
//    12'h3cc : errs =          63'b010000000000000000000000000000100000000000000000000000000000000; // D (0x2000000100000000) 
//    12'hfcc : errs =          63'b100000000000000000000000000000100000000000000000000000000000000; // D (0x4000000100000000) 
    12'haa1 : errs =          63'b000000000000000000000000000001000000000000000000000000000000001; // D (0x0000000200000001) 
    12'h5ea : errs =          63'b000000000000000000000000000001000000000000000000000000000000010; // D (0x0000000200000002) 
    12'he45 : errs =          63'b000000000000000000000000000001000000000000000000000000000000100; // D (0x0000000200000004) 
    12'hc22 : errs =          63'b000000000000000000000000000001000000000000000000000000000001000; // D (0x0000000200000008) 
    12'h8ec : errs =          63'b000000000000000000000000000001000000000000000000000000000010000; // D (0x0000000200000010) 
    12'h170 : errs =          63'b000000000000000000000000000001000000000000000000000000000100000; // D (0x0000000200000020) 
    12'h771 : errs =          63'b000000000000000000000000000001000000000000000000000000001000000; // D (0x0000000200000040) 
    12'hb73 : errs =          63'b000000000000000000000000000001000000000000000000000000010000000; // D (0x0000000200000080) 
    12'h64e : errs =          63'b000000000000000000000000000001000000000000000000000000100000000; // D (0x0000000200000100) 
    12'h90d : errs =          63'b000000000000000000000000000001000000000000000000000001000000000; // D (0x0000000200000200) 
    12'h2b2 : errs =          63'b000000000000000000000000000001000000000000000000000010000000000; // D (0x0000000200000400) 
    12'h0f5 : errs =          63'b000000000000000000000000000001000000000000000000000100000000000; // D (0x0000000200000800) 
    12'h47b : errs =          63'b000000000000000000000000000001000000000000000000001000000000000; // D (0x0000000200001000) 
    12'hd67 : errs =          63'b000000000000000000000000000001000000000000000000010000000000000; // D (0x0000000200002000) 
    12'ha66 : errs =          63'b000000000000000000000000000001000000000000000000100000000000000; // D (0x0000000200004000) 
    12'h464 : errs =          63'b000000000000000000000000000001000000000000000001000000000000000; // D (0x0000000200008000) 
    12'hd59 : errs =          63'b000000000000000000000000000001000000000000000010000000000000000; // D (0x0000000200010000) 
    12'ha1a : errs =          63'b000000000000000000000000000001000000000000000100000000000000000; // D (0x0000000200020000) 
    12'h49c : errs =          63'b000000000000000000000000000001000000000000001000000000000000000; // D (0x0000000200040000) 
    12'hca9 : errs =          63'b000000000000000000000000000001000000000000010000000000000000000; // D (0x0000000200080000) 
    12'h9fa : errs =          63'b000000000000000000000000000001000000000000100000000000000000000; // D (0x0000000200100000) 
    12'h35c : errs =          63'b000000000000000000000000000001000000000001000000000000000000000; // D (0x0000000200200000) 
    12'h329 : errs =          63'b000000000000000000000000000001000000000010000000000000000000000; // D (0x0000000200400000) 
    12'h3c3 : errs =          63'b000000000000000000000000000001000000000100000000000000000000000; // D (0x0000000200800000) 
    12'h217 : errs =          63'b000000000000000000000000000001000000001000000000000000000000000; // D (0x0000000201000000) 
    12'h1bf : errs =          63'b000000000000000000000000000001000000010000000000000000000000000; // D (0x0000000202000000) 
    12'h6ef : errs =          63'b000000000000000000000000000001000000100000000000000000000000000; // D (0x0000000204000000) 
    12'h84f : errs =          63'b000000000000000000000000000001000001000000000000000000000000000; // D (0x0000000208000000) 
    12'h036 : errs =          63'b000000000000000000000000000001000010000000000000000000000000000; // D (0x0000000210000000) 
    12'h5fd : errs =          63'b000000000000000000000000000001000100000000000000000000000000000; // D (0x0000000220000000) 
    12'he6b : errs =          63'b000000000000000000000000000001001000000000000000000000000000000; // D (0x0000000240000000) 
    12'hc7e : errs =          63'b000000000000000000000000000001010000000000000000000000000000000; // D (0x0000000280000000) 
    12'h854 : errs =          63'b000000000000000000000000000001100000000000000000000000000000000; // D (0x0000000300000000) 
    12'hf98 : errs =          63'b000000000000000000000000000001000000000000000000000000000000000; // S (0x0000000200000000) 
//    12'h591 : errs =          63'b000000000000000000000000000011000000000000000000000000000000000; // D (0x0000000600000000) 
//    12'heb3 : errs =          63'b000000000000000000000000000101000000000000000000000000000000000; // D (0x0000000a00000000) 
//    12'hdce : errs =          63'b000000000000000000000000001001000000000000000000000000000000000; // D (0x0000001200000000) 
//    12'hb34 : errs =          63'b000000000000000000000000010001000000000000000000000000000000000; // D (0x0000002200000000) 
//    12'h6c0 : errs =          63'b000000000000000000000000100001000000000000000000000000000000000; // D (0x0000004200000000) 
//    12'h811 : errs =          63'b000000000000000000000001000001000000000000000000000000000000000; // D (0x0000008200000000) 
//    12'h08a : errs =          63'b000000000000000000000010000001000000000000000000000000000000000; // D (0x0000010200000000) 
//    12'h485 : errs =          63'b000000000000000000000100000001000000000000000000000000000000000; // D (0x0000020200000000) 
//    12'hc9b : errs =          63'b000000000000000000001000000001000000000000000000000000000000000; // D (0x0000040200000000) 
//    12'h99e : errs =          63'b000000000000000000010000000001000000000000000000000000000000000; // D (0x0000080200000000) 
//    12'h394 : errs =          63'b000000000000000000100000000001000000000000000000000000000000000; // D (0x0000100200000000) 
//    12'h2b9 : errs =          63'b000000000000000001000000000001000000000000000000000000000000000; // D (0x0000200200000000) 
//    12'h0e3 : errs =          63'b000000000000000010000000000001000000000000000000000000000000000; // D (0x0000400200000000) 
//    12'h457 : errs =          63'b000000000000000100000000000001000000000000000000000000000000000; // D (0x0000800200000000) 
//    12'hd3f : errs =          63'b000000000000001000000000000001000000000000000000000000000000000; // D (0x0001000200000000) 
//    12'had6 : errs =          63'b000000000000010000000000000001000000000000000000000000000000000; // D (0x0002000200000000) 
//    12'h504 : errs =          63'b000000000000100000000000000001000000000000000000000000000000000; // D (0x0004000200000000) 
//    12'hf99 : errs =          63'b000000000001000000000000000001000000000000000000000000000000000; // D (0x0008000200000000) 
//    12'hf9a : errs =          63'b000000000010000000000000000001000000000000000000000000000000000; // D (0x0010000200000000) 
//    12'hf9c : errs =          63'b000000000100000000000000000001000000000000000000000000000000000; // D (0x0020000200000000) 
//    12'hf90 : errs =          63'b000000001000000000000000000001000000000000000000000000000000000; // D (0x0040000200000000) 
//    12'hf88 : errs =          63'b000000010000000000000000000001000000000000000000000000000000000; // D (0x0080000200000000) 
//    12'hfb8 : errs =          63'b000000100000000000000000000001000000000000000000000000000000000; // D (0x0100000200000000) 
//    12'hfd8 : errs =          63'b000001000000000000000000000001000000000000000000000000000000000; // D (0x0200000200000000) 
//    12'hf18 : errs =          63'b000010000000000000000000000001000000000000000000000000000000000; // D (0x0400000200000000) 
//    12'he98 : errs =          63'b000100000000000000000000000001000000000000000000000000000000000; // D (0x0800000200000000) 
//    12'hd98 : errs =          63'b001000000000000000000000000001000000000000000000000000000000000; // D (0x1000000200000000) 
//    12'hb98 : errs =          63'b010000000000000000000000000001000000000000000000000000000000000; // D (0x2000000200000000) 
//    12'h798 : errs =          63'b100000000000000000000000000001000000000000000000000000000000000; // D (0x4000000200000000) 
    12'hf30 : errs =          63'b000000000000000000000000000010000000000000000000000000000000001; // D (0x0000000400000001) 
    12'h07b : errs =          63'b000000000000000000000000000010000000000000000000000000000000010; // D (0x0000000400000002) 
    12'hbd4 : errs =          63'b000000000000000000000000000010000000000000000000000000000000100; // D (0x0000000400000004) 
    12'h9b3 : errs =          63'b000000000000000000000000000010000000000000000000000000000001000; // D (0x0000000400000008) 
    12'hd7d : errs =          63'b000000000000000000000000000010000000000000000000000000000010000; // D (0x0000000400000010) 
    12'h4e1 : errs =          63'b000000000000000000000000000010000000000000000000000000000100000; // D (0x0000000400000020) 
    12'h2e0 : errs =          63'b000000000000000000000000000010000000000000000000000000001000000; // D (0x0000000400000040) 
    12'hee2 : errs =          63'b000000000000000000000000000010000000000000000000000000010000000; // D (0x0000000400000080) 
    12'h3df : errs =          63'b000000000000000000000000000010000000000000000000000000100000000; // D (0x0000000400000100) 
    12'hc9c : errs =          63'b000000000000000000000000000010000000000000000000000001000000000; // D (0x0000000400000200) 
    12'h723 : errs =          63'b000000000000000000000000000010000000000000000000000010000000000; // D (0x0000000400000400) 
    12'h564 : errs =          63'b000000000000000000000000000010000000000000000000000100000000000; // D (0x0000000400000800) 
    12'h1ea : errs =          63'b000000000000000000000000000010000000000000000000001000000000000; // D (0x0000000400001000) 
    12'h8f6 : errs =          63'b000000000000000000000000000010000000000000000000010000000000000; // D (0x0000000400002000) 
    12'hff7 : errs =          63'b000000000000000000000000000010000000000000000000100000000000000; // D (0x0000000400004000) 
    12'h1f5 : errs =          63'b000000000000000000000000000010000000000000000001000000000000000; // D (0x0000000400008000) 
    12'h8c8 : errs =          63'b000000000000000000000000000010000000000000000010000000000000000; // D (0x0000000400010000) 
    12'hf8b : errs =          63'b000000000000000000000000000010000000000000000100000000000000000; // D (0x0000000400020000) 
    12'h10d : errs =          63'b000000000000000000000000000010000000000000001000000000000000000; // D (0x0000000400040000) 
    12'h938 : errs =          63'b000000000000000000000000000010000000000000010000000000000000000; // D (0x0000000400080000) 
    12'hc6b : errs =          63'b000000000000000000000000000010000000000000100000000000000000000; // D (0x0000000400100000) 
    12'h6cd : errs =          63'b000000000000000000000000000010000000000001000000000000000000000; // D (0x0000000400200000) 
    12'h6b8 : errs =          63'b000000000000000000000000000010000000000010000000000000000000000; // D (0x0000000400400000) 
    12'h652 : errs =          63'b000000000000000000000000000010000000000100000000000000000000000; // D (0x0000000400800000) 
    12'h786 : errs =          63'b000000000000000000000000000010000000001000000000000000000000000; // D (0x0000000401000000) 
    12'h42e : errs =          63'b000000000000000000000000000010000000010000000000000000000000000; // D (0x0000000402000000) 
    12'h37e : errs =          63'b000000000000000000000000000010000000100000000000000000000000000; // D (0x0000000404000000) 
    12'hdde : errs =          63'b000000000000000000000000000010000001000000000000000000000000000; // D (0x0000000408000000) 
    12'h5a7 : errs =          63'b000000000000000000000000000010000010000000000000000000000000000; // D (0x0000000410000000) 
    12'h06c : errs =          63'b000000000000000000000000000010000100000000000000000000000000000; // D (0x0000000420000000) 
    12'hbfa : errs =          63'b000000000000000000000000000010001000000000000000000000000000000; // D (0x0000000440000000) 
    12'h9ef : errs =          63'b000000000000000000000000000010010000000000000000000000000000000; // D (0x0000000480000000) 
    12'hdc5 : errs =          63'b000000000000000000000000000010100000000000000000000000000000000; // D (0x0000000500000000) 
    12'h591 : errs =          63'b000000000000000000000000000011000000000000000000000000000000000; // D (0x0000000600000000) 
    12'ha09 : errs =          63'b000000000000000000000000000010000000000000000000000000000000000; // S (0x0000000400000000) 
//    12'hb22 : errs =          63'b000000000000000000000000000110000000000000000000000000000000000; // D (0x0000000c00000000) 
//    12'h85f : errs =          63'b000000000000000000000000001010000000000000000000000000000000000; // D (0x0000001400000000) 
//    12'hea5 : errs =          63'b000000000000000000000000010010000000000000000000000000000000000; // D (0x0000002400000000) 
//    12'h351 : errs =          63'b000000000000000000000000100010000000000000000000000000000000000; // D (0x0000004400000000) 
//    12'hd80 : errs =          63'b000000000000000000000001000010000000000000000000000000000000000; // D (0x0000008400000000) 
//    12'h51b : errs =          63'b000000000000000000000010000010000000000000000000000000000000000; // D (0x0000010400000000) 
//    12'h114 : errs =          63'b000000000000000000000100000010000000000000000000000000000000000; // D (0x0000020400000000) 
//    12'h90a : errs =          63'b000000000000000000001000000010000000000000000000000000000000000; // D (0x0000040400000000) 
//    12'hc0f : errs =          63'b000000000000000000010000000010000000000000000000000000000000000; // D (0x0000080400000000) 
//    12'h605 : errs =          63'b000000000000000000100000000010000000000000000000000000000000000; // D (0x0000100400000000) 
//    12'h728 : errs =          63'b000000000000000001000000000010000000000000000000000000000000000; // D (0x0000200400000000) 
//    12'h572 : errs =          63'b000000000000000010000000000010000000000000000000000000000000000; // D (0x0000400400000000) 
//    12'h1c6 : errs =          63'b000000000000000100000000000010000000000000000000000000000000000; // D (0x0000800400000000) 
//    12'h8ae : errs =          63'b000000000000001000000000000010000000000000000000000000000000000; // D (0x0001000400000000) 
//    12'hf47 : errs =          63'b000000000000010000000000000010000000000000000000000000000000000; // D (0x0002000400000000) 
//    12'h095 : errs =          63'b000000000000100000000000000010000000000000000000000000000000000; // D (0x0004000400000000) 
//    12'ha08 : errs =          63'b000000000001000000000000000010000000000000000000000000000000000; // D (0x0008000400000000) 
//    12'ha0b : errs =          63'b000000000010000000000000000010000000000000000000000000000000000; // D (0x0010000400000000) 
//    12'ha0d : errs =          63'b000000000100000000000000000010000000000000000000000000000000000; // D (0x0020000400000000) 
//    12'ha01 : errs =          63'b000000001000000000000000000010000000000000000000000000000000000; // D (0x0040000400000000) 
//    12'ha19 : errs =          63'b000000010000000000000000000010000000000000000000000000000000000; // D (0x0080000400000000) 
//    12'ha29 : errs =          63'b000000100000000000000000000010000000000000000000000000000000000; // D (0x0100000400000000) 
//    12'ha49 : errs =          63'b000001000000000000000000000010000000000000000000000000000000000; // D (0x0200000400000000) 
//    12'ha89 : errs =          63'b000010000000000000000000000010000000000000000000000000000000000; // D (0x0400000400000000) 
//    12'hb09 : errs =          63'b000100000000000000000000000010000000000000000000000000000000000; // D (0x0800000400000000) 
//    12'h809 : errs =          63'b001000000000000000000000000010000000000000000000000000000000000; // D (0x1000000400000000) 
//    12'he09 : errs =          63'b010000000000000000000000000010000000000000000000000000000000000; // D (0x2000000400000000) 
//    12'h209 : errs =          63'b100000000000000000000000000010000000000000000000000000000000000; // D (0x4000000400000000) 
    12'h412 : errs =          63'b000000000000000000000000000100000000000000000000000000000000001; // D (0x0000000800000001) 
    12'hb59 : errs =          63'b000000000000000000000000000100000000000000000000000000000000010; // D (0x0000000800000002) 
    12'h0f6 : errs =          63'b000000000000000000000000000100000000000000000000000000000000100; // D (0x0000000800000004) 
    12'h291 : errs =          63'b000000000000000000000000000100000000000000000000000000000001000; // D (0x0000000800000008) 
    12'h65f : errs =          63'b000000000000000000000000000100000000000000000000000000000010000; // D (0x0000000800000010) 
    12'hfc3 : errs =          63'b000000000000000000000000000100000000000000000000000000000100000; // D (0x0000000800000020) 
    12'h9c2 : errs =          63'b000000000000000000000000000100000000000000000000000000001000000; // D (0x0000000800000040) 
    12'h5c0 : errs =          63'b000000000000000000000000000100000000000000000000000000010000000; // D (0x0000000800000080) 
    12'h8fd : errs =          63'b000000000000000000000000000100000000000000000000000000100000000; // D (0x0000000800000100) 
    12'h7be : errs =          63'b000000000000000000000000000100000000000000000000000001000000000; // D (0x0000000800000200) 
    12'hc01 : errs =          63'b000000000000000000000000000100000000000000000000000010000000000; // D (0x0000000800000400) 
    12'he46 : errs =          63'b000000000000000000000000000100000000000000000000000100000000000; // D (0x0000000800000800) 
    12'hac8 : errs =          63'b000000000000000000000000000100000000000000000000001000000000000; // D (0x0000000800001000) 
    12'h3d4 : errs =          63'b000000000000000000000000000100000000000000000000010000000000000; // D (0x0000000800002000) 
    12'h4d5 : errs =          63'b000000000000000000000000000100000000000000000000100000000000000; // D (0x0000000800004000) 
    12'had7 : errs =          63'b000000000000000000000000000100000000000000000001000000000000000; // D (0x0000000800008000) 
    12'h3ea : errs =          63'b000000000000000000000000000100000000000000000010000000000000000; // D (0x0000000800010000) 
    12'h4a9 : errs =          63'b000000000000000000000000000100000000000000000100000000000000000; // D (0x0000000800020000) 
    12'ha2f : errs =          63'b000000000000000000000000000100000000000000001000000000000000000; // D (0x0000000800040000) 
    12'h21a : errs =          63'b000000000000000000000000000100000000000000010000000000000000000; // D (0x0000000800080000) 
    12'h749 : errs =          63'b000000000000000000000000000100000000000000100000000000000000000; // D (0x0000000800100000) 
    12'hdef : errs =          63'b000000000000000000000000000100000000000001000000000000000000000; // D (0x0000000800200000) 
    12'hd9a : errs =          63'b000000000000000000000000000100000000000010000000000000000000000; // D (0x0000000800400000) 
    12'hd70 : errs =          63'b000000000000000000000000000100000000000100000000000000000000000; // D (0x0000000800800000) 
    12'hca4 : errs =          63'b000000000000000000000000000100000000001000000000000000000000000; // D (0x0000000801000000) 
    12'hf0c : errs =          63'b000000000000000000000000000100000000010000000000000000000000000; // D (0x0000000802000000) 
    12'h85c : errs =          63'b000000000000000000000000000100000000100000000000000000000000000; // D (0x0000000804000000) 
    12'h6fc : errs =          63'b000000000000000000000000000100000001000000000000000000000000000; // D (0x0000000808000000) 
    12'he85 : errs =          63'b000000000000000000000000000100000010000000000000000000000000000; // D (0x0000000810000000) 
    12'hb4e : errs =          63'b000000000000000000000000000100000100000000000000000000000000000; // D (0x0000000820000000) 
    12'h0d8 : errs =          63'b000000000000000000000000000100001000000000000000000000000000000; // D (0x0000000840000000) 
    12'h2cd : errs =          63'b000000000000000000000000000100010000000000000000000000000000000; // D (0x0000000880000000) 
    12'h6e7 : errs =          63'b000000000000000000000000000100100000000000000000000000000000000; // D (0x0000000900000000) 
    12'heb3 : errs =          63'b000000000000000000000000000101000000000000000000000000000000000; // D (0x0000000a00000000) 
    12'hb22 : errs =          63'b000000000000000000000000000110000000000000000000000000000000000; // D (0x0000000c00000000) 
    12'h12b : errs =          63'b000000000000000000000000000100000000000000000000000000000000000; // S (0x0000000800000000) 
//    12'h37d : errs =          63'b000000000000000000000000001100000000000000000000000000000000000; // D (0x0000001800000000) 
//    12'h587 : errs =          63'b000000000000000000000000010100000000000000000000000000000000000; // D (0x0000002800000000) 
//    12'h873 : errs =          63'b000000000000000000000000100100000000000000000000000000000000000; // D (0x0000004800000000) 
//    12'h6a2 : errs =          63'b000000000000000000000001000100000000000000000000000000000000000; // D (0x0000008800000000) 
//    12'he39 : errs =          63'b000000000000000000000010000100000000000000000000000000000000000; // D (0x0000010800000000) 
//    12'ha36 : errs =          63'b000000000000000000000100000100000000000000000000000000000000000; // D (0x0000020800000000) 
//    12'h228 : errs =          63'b000000000000000000001000000100000000000000000000000000000000000; // D (0x0000040800000000) 
//    12'h72d : errs =          63'b000000000000000000010000000100000000000000000000000000000000000; // D (0x0000080800000000) 
//    12'hd27 : errs =          63'b000000000000000000100000000100000000000000000000000000000000000; // D (0x0000100800000000) 
//    12'hc0a : errs =          63'b000000000000000001000000000100000000000000000000000000000000000; // D (0x0000200800000000) 
//    12'he50 : errs =          63'b000000000000000010000000000100000000000000000000000000000000000; // D (0x0000400800000000) 
//    12'hae4 : errs =          63'b000000000000000100000000000100000000000000000000000000000000000; // D (0x0000800800000000) 
//    12'h38c : errs =          63'b000000000000001000000000000100000000000000000000000000000000000; // D (0x0001000800000000) 
//    12'h465 : errs =          63'b000000000000010000000000000100000000000000000000000000000000000; // D (0x0002000800000000) 
//    12'hbb7 : errs =          63'b000000000000100000000000000100000000000000000000000000000000000; // D (0x0004000800000000) 
//    12'h12a : errs =          63'b000000000001000000000000000100000000000000000000000000000000000; // D (0x0008000800000000) 
//    12'h129 : errs =          63'b000000000010000000000000000100000000000000000000000000000000000; // D (0x0010000800000000) 
//    12'h12f : errs =          63'b000000000100000000000000000100000000000000000000000000000000000; // D (0x0020000800000000) 
//    12'h123 : errs =          63'b000000001000000000000000000100000000000000000000000000000000000; // D (0x0040000800000000) 
//    12'h13b : errs =          63'b000000010000000000000000000100000000000000000000000000000000000; // D (0x0080000800000000) 
//    12'h10b : errs =          63'b000000100000000000000000000100000000000000000000000000000000000; // D (0x0100000800000000) 
//    12'h16b : errs =          63'b000001000000000000000000000100000000000000000000000000000000000; // D (0x0200000800000000) 
//    12'h1ab : errs =          63'b000010000000000000000000000100000000000000000000000000000000000; // D (0x0400000800000000) 
//    12'h02b : errs =          63'b000100000000000000000000000100000000000000000000000000000000000; // D (0x0800000800000000) 
//    12'h32b : errs =          63'b001000000000000000000000000100000000000000000000000000000000000; // D (0x1000000800000000) 
//    12'h52b : errs =          63'b010000000000000000000000000100000000000000000000000000000000000; // D (0x2000000800000000) 
//    12'h92b : errs =          63'b100000000000000000000000000100000000000000000000000000000000000; // D (0x4000000800000000) 
    12'h76f : errs =          63'b000000000000000000000000001000000000000000000000000000000000001; // D (0x0000001000000001) 
    12'h824 : errs =          63'b000000000000000000000000001000000000000000000000000000000000010; // D (0x0000001000000002) 
    12'h38b : errs =          63'b000000000000000000000000001000000000000000000000000000000000100; // D (0x0000001000000004) 
    12'h1ec : errs =          63'b000000000000000000000000001000000000000000000000000000000001000; // D (0x0000001000000008) 
    12'h522 : errs =          63'b000000000000000000000000001000000000000000000000000000000010000; // D (0x0000001000000010) 
    12'hcbe : errs =          63'b000000000000000000000000001000000000000000000000000000000100000; // D (0x0000001000000020) 
    12'habf : errs =          63'b000000000000000000000000001000000000000000000000000000001000000; // D (0x0000001000000040) 
    12'h6bd : errs =          63'b000000000000000000000000001000000000000000000000000000010000000; // D (0x0000001000000080) 
    12'hb80 : errs =          63'b000000000000000000000000001000000000000000000000000000100000000; // D (0x0000001000000100) 
    12'h4c3 : errs =          63'b000000000000000000000000001000000000000000000000000001000000000; // D (0x0000001000000200) 
    12'hf7c : errs =          63'b000000000000000000000000001000000000000000000000000010000000000; // D (0x0000001000000400) 
    12'hd3b : errs =          63'b000000000000000000000000001000000000000000000000000100000000000; // D (0x0000001000000800) 
    12'h9b5 : errs =          63'b000000000000000000000000001000000000000000000000001000000000000; // D (0x0000001000001000) 
    12'h0a9 : errs =          63'b000000000000000000000000001000000000000000000000010000000000000; // D (0x0000001000002000) 
    12'h7a8 : errs =          63'b000000000000000000000000001000000000000000000000100000000000000; // D (0x0000001000004000) 
    12'h9aa : errs =          63'b000000000000000000000000001000000000000000000001000000000000000; // D (0x0000001000008000) 
    12'h097 : errs =          63'b000000000000000000000000001000000000000000000010000000000000000; // D (0x0000001000010000) 
    12'h7d4 : errs =          63'b000000000000000000000000001000000000000000000100000000000000000; // D (0x0000001000020000) 
    12'h952 : errs =          63'b000000000000000000000000001000000000000000001000000000000000000; // D (0x0000001000040000) 
    12'h167 : errs =          63'b000000000000000000000000001000000000000000010000000000000000000; // D (0x0000001000080000) 
    12'h434 : errs =          63'b000000000000000000000000001000000000000000100000000000000000000; // D (0x0000001000100000) 
    12'he92 : errs =          63'b000000000000000000000000001000000000000001000000000000000000000; // D (0x0000001000200000) 
    12'hee7 : errs =          63'b000000000000000000000000001000000000000010000000000000000000000; // D (0x0000001000400000) 
    12'he0d : errs =          63'b000000000000000000000000001000000000000100000000000000000000000; // D (0x0000001000800000) 
    12'hfd9 : errs =          63'b000000000000000000000000001000000000001000000000000000000000000; // D (0x0000001001000000) 
    12'hc71 : errs =          63'b000000000000000000000000001000000000010000000000000000000000000; // D (0x0000001002000000) 
    12'hb21 : errs =          63'b000000000000000000000000001000000000100000000000000000000000000; // D (0x0000001004000000) 
    12'h581 : errs =          63'b000000000000000000000000001000000001000000000000000000000000000; // D (0x0000001008000000) 
    12'hdf8 : errs =          63'b000000000000000000000000001000000010000000000000000000000000000; // D (0x0000001010000000) 
    12'h833 : errs =          63'b000000000000000000000000001000000100000000000000000000000000000; // D (0x0000001020000000) 
    12'h3a5 : errs =          63'b000000000000000000000000001000001000000000000000000000000000000; // D (0x0000001040000000) 
    12'h1b0 : errs =          63'b000000000000000000000000001000010000000000000000000000000000000; // D (0x0000001080000000) 
    12'h59a : errs =          63'b000000000000000000000000001000100000000000000000000000000000000; // D (0x0000001100000000) 
    12'hdce : errs =          63'b000000000000000000000000001001000000000000000000000000000000000; // D (0x0000001200000000) 
    12'h85f : errs =          63'b000000000000000000000000001010000000000000000000000000000000000; // D (0x0000001400000000) 
    12'h37d : errs =          63'b000000000000000000000000001100000000000000000000000000000000000; // D (0x0000001800000000) 
    12'h256 : errs =          63'b000000000000000000000000001000000000000000000000000000000000000; // S (0x0000001000000000) 
//    12'h6fa : errs =          63'b000000000000000000000000011000000000000000000000000000000000000; // D (0x0000003000000000) 
//    12'hb0e : errs =          63'b000000000000000000000000101000000000000000000000000000000000000; // D (0x0000005000000000) 
//    12'h5df : errs =          63'b000000000000000000000001001000000000000000000000000000000000000; // D (0x0000009000000000) 
//    12'hd44 : errs =          63'b000000000000000000000010001000000000000000000000000000000000000; // D (0x0000011000000000) 
//    12'h94b : errs =          63'b000000000000000000000100001000000000000000000000000000000000000; // D (0x0000021000000000) 
//    12'h155 : errs =          63'b000000000000000000001000001000000000000000000000000000000000000; // D (0x0000041000000000) 
//    12'h450 : errs =          63'b000000000000000000010000001000000000000000000000000000000000000; // D (0x0000081000000000) 
//    12'he5a : errs =          63'b000000000000000000100000001000000000000000000000000000000000000; // D (0x0000101000000000) 
//    12'hf77 : errs =          63'b000000000000000001000000001000000000000000000000000000000000000; // D (0x0000201000000000) 
//    12'hd2d : errs =          63'b000000000000000010000000001000000000000000000000000000000000000; // D (0x0000401000000000) 
//    12'h999 : errs =          63'b000000000000000100000000001000000000000000000000000000000000000; // D (0x0000801000000000) 
//    12'h0f1 : errs =          63'b000000000000001000000000001000000000000000000000000000000000000; // D (0x0001001000000000) 
//    12'h718 : errs =          63'b000000000000010000000000001000000000000000000000000000000000000; // D (0x0002001000000000) 
//    12'h8ca : errs =          63'b000000000000100000000000001000000000000000000000000000000000000; // D (0x0004001000000000) 
//    12'h257 : errs =          63'b000000000001000000000000001000000000000000000000000000000000000; // D (0x0008001000000000) 
//    12'h254 : errs =          63'b000000000010000000000000001000000000000000000000000000000000000; // D (0x0010001000000000) 
//    12'h252 : errs =          63'b000000000100000000000000001000000000000000000000000000000000000; // D (0x0020001000000000) 
//    12'h25e : errs =          63'b000000001000000000000000001000000000000000000000000000000000000; // D (0x0040001000000000) 
//    12'h246 : errs =          63'b000000010000000000000000001000000000000000000000000000000000000; // D (0x0080001000000000) 
//    12'h276 : errs =          63'b000000100000000000000000001000000000000000000000000000000000000; // D (0x0100001000000000) 
//    12'h216 : errs =          63'b000001000000000000000000001000000000000000000000000000000000000; // D (0x0200001000000000) 
//    12'h2d6 : errs =          63'b000010000000000000000000001000000000000000000000000000000000000; // D (0x0400001000000000) 
//    12'h356 : errs =          63'b000100000000000000000000001000000000000000000000000000000000000; // D (0x0800001000000000) 
//    12'h056 : errs =          63'b001000000000000000000000001000000000000000000000000000000000000; // D (0x1000001000000000) 
//    12'h656 : errs =          63'b010000000000000000000000001000000000000000000000000000000000000; // D (0x2000001000000000) 
//    12'ha56 : errs =          63'b100000000000000000000000001000000000000000000000000000000000000; // D (0x4000001000000000) 
    12'h195 : errs =          63'b000000000000000000000000010000000000000000000000000000000000001; // D (0x0000002000000001) 
    12'hede : errs =          63'b000000000000000000000000010000000000000000000000000000000000010; // D (0x0000002000000002) 
    12'h571 : errs =          63'b000000000000000000000000010000000000000000000000000000000000100; // D (0x0000002000000004) 
    12'h716 : errs =          63'b000000000000000000000000010000000000000000000000000000000001000; // D (0x0000002000000008) 
    12'h3d8 : errs =          63'b000000000000000000000000010000000000000000000000000000000010000; // D (0x0000002000000010) 
    12'ha44 : errs =          63'b000000000000000000000000010000000000000000000000000000000100000; // D (0x0000002000000020) 
    12'hc45 : errs =          63'b000000000000000000000000010000000000000000000000000000001000000; // D (0x0000002000000040) 
    12'h047 : errs =          63'b000000000000000000000000010000000000000000000000000000010000000; // D (0x0000002000000080) 
    12'hd7a : errs =          63'b000000000000000000000000010000000000000000000000000000100000000; // D (0x0000002000000100) 
    12'h239 : errs =          63'b000000000000000000000000010000000000000000000000000001000000000; // D (0x0000002000000200) 
    12'h986 : errs =          63'b000000000000000000000000010000000000000000000000000010000000000; // D (0x0000002000000400) 
    12'hbc1 : errs =          63'b000000000000000000000000010000000000000000000000000100000000000; // D (0x0000002000000800) 
    12'hf4f : errs =          63'b000000000000000000000000010000000000000000000000001000000000000; // D (0x0000002000001000) 
    12'h653 : errs =          63'b000000000000000000000000010000000000000000000000010000000000000; // D (0x0000002000002000) 
    12'h152 : errs =          63'b000000000000000000000000010000000000000000000000100000000000000; // D (0x0000002000004000) 
    12'hf50 : errs =          63'b000000000000000000000000010000000000000000000001000000000000000; // D (0x0000002000008000) 
    12'h66d : errs =          63'b000000000000000000000000010000000000000000000010000000000000000; // D (0x0000002000010000) 
    12'h12e : errs =          63'b000000000000000000000000010000000000000000000100000000000000000; // D (0x0000002000020000) 
    12'hfa8 : errs =          63'b000000000000000000000000010000000000000000001000000000000000000; // D (0x0000002000040000) 
    12'h79d : errs =          63'b000000000000000000000000010000000000000000010000000000000000000; // D (0x0000002000080000) 
    12'h2ce : errs =          63'b000000000000000000000000010000000000000000100000000000000000000; // D (0x0000002000100000) 
    12'h868 : errs =          63'b000000000000000000000000010000000000000001000000000000000000000; // D (0x0000002000200000) 
    12'h81d : errs =          63'b000000000000000000000000010000000000000010000000000000000000000; // D (0x0000002000400000) 
    12'h8f7 : errs =          63'b000000000000000000000000010000000000000100000000000000000000000; // D (0x0000002000800000) 
    12'h923 : errs =          63'b000000000000000000000000010000000000001000000000000000000000000; // D (0x0000002001000000) 
    12'ha8b : errs =          63'b000000000000000000000000010000000000010000000000000000000000000; // D (0x0000002002000000) 
    12'hddb : errs =          63'b000000000000000000000000010000000000100000000000000000000000000; // D (0x0000002004000000) 
    12'h37b : errs =          63'b000000000000000000000000010000000001000000000000000000000000000; // D (0x0000002008000000) 
    12'hb02 : errs =          63'b000000000000000000000000010000000010000000000000000000000000000; // D (0x0000002010000000) 
    12'hec9 : errs =          63'b000000000000000000000000010000000100000000000000000000000000000; // D (0x0000002020000000) 
    12'h55f : errs =          63'b000000000000000000000000010000001000000000000000000000000000000; // D (0x0000002040000000) 
    12'h74a : errs =          63'b000000000000000000000000010000010000000000000000000000000000000; // D (0x0000002080000000) 
    12'h360 : errs =          63'b000000000000000000000000010000100000000000000000000000000000000; // D (0x0000002100000000) 
    12'hb34 : errs =          63'b000000000000000000000000010001000000000000000000000000000000000; // D (0x0000002200000000) 
    12'hea5 : errs =          63'b000000000000000000000000010010000000000000000000000000000000000; // D (0x0000002400000000) 
    12'h587 : errs =          63'b000000000000000000000000010100000000000000000000000000000000000; // D (0x0000002800000000) 
    12'h6fa : errs =          63'b000000000000000000000000011000000000000000000000000000000000000; // D (0x0000003000000000) 
    12'h4ac : errs =          63'b000000000000000000000000010000000000000000000000000000000000000; // S (0x0000002000000000) 
//    12'hdf4 : errs =          63'b000000000000000000000000110000000000000000000000000000000000000; // D (0x0000006000000000) 
//    12'h325 : errs =          63'b000000000000000000000001010000000000000000000000000000000000000; // D (0x000000a000000000) 
//    12'hbbe : errs =          63'b000000000000000000000010010000000000000000000000000000000000000; // D (0x0000012000000000) 
//    12'hfb1 : errs =          63'b000000000000000000000100010000000000000000000000000000000000000; // D (0x0000022000000000) 
//    12'h7af : errs =          63'b000000000000000000001000010000000000000000000000000000000000000; // D (0x0000042000000000) 
//    12'h2aa : errs =          63'b000000000000000000010000010000000000000000000000000000000000000; // D (0x0000082000000000) 
//    12'h8a0 : errs =          63'b000000000000000000100000010000000000000000000000000000000000000; // D (0x0000102000000000) 
//    12'h98d : errs =          63'b000000000000000001000000010000000000000000000000000000000000000; // D (0x0000202000000000) 
//    12'hbd7 : errs =          63'b000000000000000010000000010000000000000000000000000000000000000; // D (0x0000402000000000) 
//    12'hf63 : errs =          63'b000000000000000100000000010000000000000000000000000000000000000; // D (0x0000802000000000) 
//    12'h60b : errs =          63'b000000000000001000000000010000000000000000000000000000000000000; // D (0x0001002000000000) 
//    12'h1e2 : errs =          63'b000000000000010000000000010000000000000000000000000000000000000; // D (0x0002002000000000) 
//    12'he30 : errs =          63'b000000000000100000000000010000000000000000000000000000000000000; // D (0x0004002000000000) 
//    12'h4ad : errs =          63'b000000000001000000000000010000000000000000000000000000000000000; // D (0x0008002000000000) 
//    12'h4ae : errs =          63'b000000000010000000000000010000000000000000000000000000000000000; // D (0x0010002000000000) 
//    12'h4a8 : errs =          63'b000000000100000000000000010000000000000000000000000000000000000; // D (0x0020002000000000) 
//    12'h4a4 : errs =          63'b000000001000000000000000010000000000000000000000000000000000000; // D (0x0040002000000000) 
//    12'h4bc : errs =          63'b000000010000000000000000010000000000000000000000000000000000000; // D (0x0080002000000000) 
//    12'h48c : errs =          63'b000000100000000000000000010000000000000000000000000000000000000; // D (0x0100002000000000) 
//    12'h4ec : errs =          63'b000001000000000000000000010000000000000000000000000000000000000; // D (0x0200002000000000) 
//    12'h42c : errs =          63'b000010000000000000000000010000000000000000000000000000000000000; // D (0x0400002000000000) 
//    12'h5ac : errs =          63'b000100000000000000000000010000000000000000000000000000000000000; // D (0x0800002000000000) 
//    12'h6ac : errs =          63'b001000000000000000000000010000000000000000000000000000000000000; // D (0x1000002000000000) 
//    12'h0ac : errs =          63'b010000000000000000000000010000000000000000000000000000000000000; // D (0x2000002000000000) 
//    12'hcac : errs =          63'b100000000000000000000000010000000000000000000000000000000000000; // D (0x4000002000000000) 
    12'hc61 : errs =          63'b000000000000000000000000100000000000000000000000000000000000001; // D (0x0000004000000001) 
    12'h32a : errs =          63'b000000000000000000000000100000000000000000000000000000000000010; // D (0x0000004000000002) 
    12'h885 : errs =          63'b000000000000000000000000100000000000000000000000000000000000100; // D (0x0000004000000004) 
    12'hae2 : errs =          63'b000000000000000000000000100000000000000000000000000000000001000; // D (0x0000004000000008) 
    12'he2c : errs =          63'b000000000000000000000000100000000000000000000000000000000010000; // D (0x0000004000000010) 
    12'h7b0 : errs =          63'b000000000000000000000000100000000000000000000000000000000100000; // D (0x0000004000000020) 
    12'h1b1 : errs =          63'b000000000000000000000000100000000000000000000000000000001000000; // D (0x0000004000000040) 
    12'hdb3 : errs =          63'b000000000000000000000000100000000000000000000000000000010000000; // D (0x0000004000000080) 
    12'h08e : errs =          63'b000000000000000000000000100000000000000000000000000000100000000; // D (0x0000004000000100) 
    12'hfcd : errs =          63'b000000000000000000000000100000000000000000000000000001000000000; // D (0x0000004000000200) 
    12'h472 : errs =          63'b000000000000000000000000100000000000000000000000000010000000000; // D (0x0000004000000400) 
    12'h635 : errs =          63'b000000000000000000000000100000000000000000000000000100000000000; // D (0x0000004000000800) 
    12'h2bb : errs =          63'b000000000000000000000000100000000000000000000000001000000000000; // D (0x0000004000001000) 
    12'hba7 : errs =          63'b000000000000000000000000100000000000000000000000010000000000000; // D (0x0000004000002000) 
    12'hca6 : errs =          63'b000000000000000000000000100000000000000000000000100000000000000; // D (0x0000004000004000) 
    12'h2a4 : errs =          63'b000000000000000000000000100000000000000000000001000000000000000; // D (0x0000004000008000) 
    12'hb99 : errs =          63'b000000000000000000000000100000000000000000000010000000000000000; // D (0x0000004000010000) 
    12'hcda : errs =          63'b000000000000000000000000100000000000000000000100000000000000000; // D (0x0000004000020000) 
    12'h25c : errs =          63'b000000000000000000000000100000000000000000001000000000000000000; // D (0x0000004000040000) 
    12'ha69 : errs =          63'b000000000000000000000000100000000000000000010000000000000000000; // D (0x0000004000080000) 
    12'hf3a : errs =          63'b000000000000000000000000100000000000000000100000000000000000000; // D (0x0000004000100000) 
    12'h59c : errs =          63'b000000000000000000000000100000000000000001000000000000000000000; // D (0x0000004000200000) 
    12'h5e9 : errs =          63'b000000000000000000000000100000000000000010000000000000000000000; // D (0x0000004000400000) 
    12'h503 : errs =          63'b000000000000000000000000100000000000000100000000000000000000000; // D (0x0000004000800000) 
    12'h4d7 : errs =          63'b000000000000000000000000100000000000001000000000000000000000000; // D (0x0000004001000000) 
    12'h77f : errs =          63'b000000000000000000000000100000000000010000000000000000000000000; // D (0x0000004002000000) 
    12'h02f : errs =          63'b000000000000000000000000100000000000100000000000000000000000000; // D (0x0000004004000000) 
    12'he8f : errs =          63'b000000000000000000000000100000000001000000000000000000000000000; // D (0x0000004008000000) 
    12'h6f6 : errs =          63'b000000000000000000000000100000000010000000000000000000000000000; // D (0x0000004010000000) 
    12'h33d : errs =          63'b000000000000000000000000100000000100000000000000000000000000000; // D (0x0000004020000000) 
    12'h8ab : errs =          63'b000000000000000000000000100000001000000000000000000000000000000; // D (0x0000004040000000) 
    12'habe : errs =          63'b000000000000000000000000100000010000000000000000000000000000000; // D (0x0000004080000000) 
    12'he94 : errs =          63'b000000000000000000000000100000100000000000000000000000000000000; // D (0x0000004100000000) 
    12'h6c0 : errs =          63'b000000000000000000000000100001000000000000000000000000000000000; // D (0x0000004200000000) 
    12'h351 : errs =          63'b000000000000000000000000100010000000000000000000000000000000000; // D (0x0000004400000000) 
    12'h873 : errs =          63'b000000000000000000000000100100000000000000000000000000000000000; // D (0x0000004800000000) 
    12'hb0e : errs =          63'b000000000000000000000000101000000000000000000000000000000000000; // D (0x0000005000000000) 
    12'hdf4 : errs =          63'b000000000000000000000000110000000000000000000000000000000000000; // D (0x0000006000000000) 
    12'h958 : errs =          63'b000000000000000000000000100000000000000000000000000000000000000; // S (0x0000004000000000) 
//    12'hed1 : errs =          63'b000000000000000000000001100000000000000000000000000000000000000; // D (0x000000c000000000) 
//    12'h64a : errs =          63'b000000000000000000000010100000000000000000000000000000000000000; // D (0x0000014000000000) 
//    12'h245 : errs =          63'b000000000000000000000100100000000000000000000000000000000000000; // D (0x0000024000000000) 
//    12'ha5b : errs =          63'b000000000000000000001000100000000000000000000000000000000000000; // D (0x0000044000000000) 
//    12'hf5e : errs =          63'b000000000000000000010000100000000000000000000000000000000000000; // D (0x0000084000000000) 
//    12'h554 : errs =          63'b000000000000000000100000100000000000000000000000000000000000000; // D (0x0000104000000000) 
//    12'h479 : errs =          63'b000000000000000001000000100000000000000000000000000000000000000; // D (0x0000204000000000) 
//    12'h623 : errs =          63'b000000000000000010000000100000000000000000000000000000000000000; // D (0x0000404000000000) 
//    12'h297 : errs =          63'b000000000000000100000000100000000000000000000000000000000000000; // D (0x0000804000000000) 
//    12'hbff : errs =          63'b000000000000001000000000100000000000000000000000000000000000000; // D (0x0001004000000000) 
//    12'hc16 : errs =          63'b000000000000010000000000100000000000000000000000000000000000000; // D (0x0002004000000000) 
//    12'h3c4 : errs =          63'b000000000000100000000000100000000000000000000000000000000000000; // D (0x0004004000000000) 
//    12'h959 : errs =          63'b000000000001000000000000100000000000000000000000000000000000000; // D (0x0008004000000000) 
//    12'h95a : errs =          63'b000000000010000000000000100000000000000000000000000000000000000; // D (0x0010004000000000) 
//    12'h95c : errs =          63'b000000000100000000000000100000000000000000000000000000000000000; // D (0x0020004000000000) 
//    12'h950 : errs =          63'b000000001000000000000000100000000000000000000000000000000000000; // D (0x0040004000000000) 
//    12'h948 : errs =          63'b000000010000000000000000100000000000000000000000000000000000000; // D (0x0080004000000000) 
//    12'h978 : errs =          63'b000000100000000000000000100000000000000000000000000000000000000; // D (0x0100004000000000) 
//    12'h918 : errs =          63'b000001000000000000000000100000000000000000000000000000000000000; // D (0x0200004000000000) 
//    12'h9d8 : errs =          63'b000010000000000000000000100000000000000000000000000000000000000; // D (0x0400004000000000) 
//    12'h858 : errs =          63'b000100000000000000000000100000000000000000000000000000000000000; // D (0x0800004000000000) 
//    12'hb58 : errs =          63'b001000000000000000000000100000000000000000000000000000000000000; // D (0x1000004000000000) 
//    12'hd58 : errs =          63'b010000000000000000000000100000000000000000000000000000000000000; // D (0x2000004000000000) 
//    12'h158 : errs =          63'b100000000000000000000000100000000000000000000000000000000000000; // D (0x4000004000000000) 
    12'h2b0 : errs =          63'b000000000000000000000001000000000000000000000000000000000000001; // D (0x0000008000000001) 
    12'hdfb : errs =          63'b000000000000000000000001000000000000000000000000000000000000010; // D (0x0000008000000002) 
    12'h654 : errs =          63'b000000000000000000000001000000000000000000000000000000000000100; // D (0x0000008000000004) 
    12'h433 : errs =          63'b000000000000000000000001000000000000000000000000000000000001000; // D (0x0000008000000008) 
    12'h0fd : errs =          63'b000000000000000000000001000000000000000000000000000000000010000; // D (0x0000008000000010) 
    12'h961 : errs =          63'b000000000000000000000001000000000000000000000000000000000100000; // D (0x0000008000000020) 
    12'hf60 : errs =          63'b000000000000000000000001000000000000000000000000000000001000000; // D (0x0000008000000040) 
    12'h362 : errs =          63'b000000000000000000000001000000000000000000000000000000010000000; // D (0x0000008000000080) 
    12'he5f : errs =          63'b000000000000000000000001000000000000000000000000000000100000000; // D (0x0000008000000100) 
    12'h11c : errs =          63'b000000000000000000000001000000000000000000000000000001000000000; // D (0x0000008000000200) 
    12'haa3 : errs =          63'b000000000000000000000001000000000000000000000000000010000000000; // D (0x0000008000000400) 
    12'h8e4 : errs =          63'b000000000000000000000001000000000000000000000000000100000000000; // D (0x0000008000000800) 
    12'hc6a : errs =          63'b000000000000000000000001000000000000000000000000001000000000000; // D (0x0000008000001000) 
    12'h576 : errs =          63'b000000000000000000000001000000000000000000000000010000000000000; // D (0x0000008000002000) 
    12'h277 : errs =          63'b000000000000000000000001000000000000000000000000100000000000000; // D (0x0000008000004000) 
    12'hc75 : errs =          63'b000000000000000000000001000000000000000000000001000000000000000; // D (0x0000008000008000) 
    12'h548 : errs =          63'b000000000000000000000001000000000000000000000010000000000000000; // D (0x0000008000010000) 
    12'h20b : errs =          63'b000000000000000000000001000000000000000000000100000000000000000; // D (0x0000008000020000) 
    12'hc8d : errs =          63'b000000000000000000000001000000000000000000001000000000000000000; // D (0x0000008000040000) 
    12'h4b8 : errs =          63'b000000000000000000000001000000000000000000010000000000000000000; // D (0x0000008000080000) 
    12'h1eb : errs =          63'b000000000000000000000001000000000000000000100000000000000000000; // D (0x0000008000100000) 
    12'hb4d : errs =          63'b000000000000000000000001000000000000000001000000000000000000000; // D (0x0000008000200000) 
    12'hb38 : errs =          63'b000000000000000000000001000000000000000010000000000000000000000; // D (0x0000008000400000) 
    12'hbd2 : errs =          63'b000000000000000000000001000000000000000100000000000000000000000; // D (0x0000008000800000) 
    12'ha06 : errs =          63'b000000000000000000000001000000000000001000000000000000000000000; // D (0x0000008001000000) 
    12'h9ae : errs =          63'b000000000000000000000001000000000000010000000000000000000000000; // D (0x0000008002000000) 
    12'hefe : errs =          63'b000000000000000000000001000000000000100000000000000000000000000; // D (0x0000008004000000) 
    12'h05e : errs =          63'b000000000000000000000001000000000001000000000000000000000000000; // D (0x0000008008000000) 
    12'h827 : errs =          63'b000000000000000000000001000000000010000000000000000000000000000; // D (0x0000008010000000) 
    12'hdec : errs =          63'b000000000000000000000001000000000100000000000000000000000000000; // D (0x0000008020000000) 
    12'h67a : errs =          63'b000000000000000000000001000000001000000000000000000000000000000; // D (0x0000008040000000) 
    12'h46f : errs =          63'b000000000000000000000001000000010000000000000000000000000000000; // D (0x0000008080000000) 
    12'h045 : errs =          63'b000000000000000000000001000000100000000000000000000000000000000; // D (0x0000008100000000) 
    12'h811 : errs =          63'b000000000000000000000001000001000000000000000000000000000000000; // D (0x0000008200000000) 
    12'hd80 : errs =          63'b000000000000000000000001000010000000000000000000000000000000000; // D (0x0000008400000000) 
    12'h6a2 : errs =          63'b000000000000000000000001000100000000000000000000000000000000000; // D (0x0000008800000000) 
    12'h5df : errs =          63'b000000000000000000000001001000000000000000000000000000000000000; // D (0x0000009000000000) 
    12'h325 : errs =          63'b000000000000000000000001010000000000000000000000000000000000000; // D (0x000000a000000000) 
    12'hed1 : errs =          63'b000000000000000000000001100000000000000000000000000000000000000; // D (0x000000c000000000) 
    12'h789 : errs =          63'b000000000000000000000001000000000000000000000000000000000000000; // S (0x0000008000000000) 
//    12'h89b : errs =          63'b000000000000000000000011000000000000000000000000000000000000000; // D (0x0000018000000000) 
//    12'hc94 : errs =          63'b000000000000000000000101000000000000000000000000000000000000000; // D (0x0000028000000000) 
//    12'h48a : errs =          63'b000000000000000000001001000000000000000000000000000000000000000; // D (0x0000048000000000) 
//    12'h18f : errs =          63'b000000000000000000010001000000000000000000000000000000000000000; // D (0x0000088000000000) 
//    12'hb85 : errs =          63'b000000000000000000100001000000000000000000000000000000000000000; // D (0x0000108000000000) 
//    12'haa8 : errs =          63'b000000000000000001000001000000000000000000000000000000000000000; // D (0x0000208000000000) 
//    12'h8f2 : errs =          63'b000000000000000010000001000000000000000000000000000000000000000; // D (0x0000408000000000) 
//    12'hc46 : errs =          63'b000000000000000100000001000000000000000000000000000000000000000; // D (0x0000808000000000) 
//    12'h52e : errs =          63'b000000000000001000000001000000000000000000000000000000000000000; // D (0x0001008000000000) 
//    12'h2c7 : errs =          63'b000000000000010000000001000000000000000000000000000000000000000; // D (0x0002008000000000) 
//    12'hd15 : errs =          63'b000000000000100000000001000000000000000000000000000000000000000; // D (0x0004008000000000) 
//    12'h788 : errs =          63'b000000000001000000000001000000000000000000000000000000000000000; // D (0x0008008000000000) 
//    12'h78b : errs =          63'b000000000010000000000001000000000000000000000000000000000000000; // D (0x0010008000000000) 
//    12'h78d : errs =          63'b000000000100000000000001000000000000000000000000000000000000000; // D (0x0020008000000000) 
//    12'h781 : errs =          63'b000000001000000000000001000000000000000000000000000000000000000; // D (0x0040008000000000) 
//    12'h799 : errs =          63'b000000010000000000000001000000000000000000000000000000000000000; // D (0x0080008000000000) 
//    12'h7a9 : errs =          63'b000000100000000000000001000000000000000000000000000000000000000; // D (0x0100008000000000) 
//    12'h7c9 : errs =          63'b000001000000000000000001000000000000000000000000000000000000000; // D (0x0200008000000000) 
//    12'h709 : errs =          63'b000010000000000000000001000000000000000000000000000000000000000; // D (0x0400008000000000) 
//    12'h689 : errs =          63'b000100000000000000000001000000000000000000000000000000000000000; // D (0x0800008000000000) 
//    12'h589 : errs =          63'b001000000000000000000001000000000000000000000000000000000000000; // D (0x1000008000000000) 
//    12'h389 : errs =          63'b010000000000000000000001000000000000000000000000000000000000000; // D (0x2000008000000000) 
//    12'hf89 : errs =          63'b100000000000000000000001000000000000000000000000000000000000000; // D (0x4000008000000000) 
    12'ha2b : errs =          63'b000000000000000000000010000000000000000000000000000000000000001; // D (0x0000010000000001) 
    12'h560 : errs =          63'b000000000000000000000010000000000000000000000000000000000000010; // D (0x0000010000000002) 
    12'hecf : errs =          63'b000000000000000000000010000000000000000000000000000000000000100; // D (0x0000010000000004) 
    12'hca8 : errs =          63'b000000000000000000000010000000000000000000000000000000000001000; // D (0x0000010000000008) 
    12'h866 : errs =          63'b000000000000000000000010000000000000000000000000000000000010000; // D (0x0000010000000010) 
    12'h1fa : errs =          63'b000000000000000000000010000000000000000000000000000000000100000; // D (0x0000010000000020) 
    12'h7fb : errs =          63'b000000000000000000000010000000000000000000000000000000001000000; // D (0x0000010000000040) 
    12'hbf9 : errs =          63'b000000000000000000000010000000000000000000000000000000010000000; // D (0x0000010000000080) 
    12'h6c4 : errs =          63'b000000000000000000000010000000000000000000000000000000100000000; // D (0x0000010000000100) 
    12'h987 : errs =          63'b000000000000000000000010000000000000000000000000000001000000000; // D (0x0000010000000200) 
    12'h238 : errs =          63'b000000000000000000000010000000000000000000000000000010000000000; // D (0x0000010000000400) 
    12'h07f : errs =          63'b000000000000000000000010000000000000000000000000000100000000000; // D (0x0000010000000800) 
    12'h4f1 : errs =          63'b000000000000000000000010000000000000000000000000001000000000000; // D (0x0000010000001000) 
    12'hded : errs =          63'b000000000000000000000010000000000000000000000000010000000000000; // D (0x0000010000002000) 
    12'haec : errs =          63'b000000000000000000000010000000000000000000000000100000000000000; // D (0x0000010000004000) 
    12'h4ee : errs =          63'b000000000000000000000010000000000000000000000001000000000000000; // D (0x0000010000008000) 
    12'hdd3 : errs =          63'b000000000000000000000010000000000000000000000010000000000000000; // D (0x0000010000010000) 
    12'ha90 : errs =          63'b000000000000000000000010000000000000000000000100000000000000000; // D (0x0000010000020000) 
    12'h416 : errs =          63'b000000000000000000000010000000000000000000001000000000000000000; // D (0x0000010000040000) 
    12'hc23 : errs =          63'b000000000000000000000010000000000000000000010000000000000000000; // D (0x0000010000080000) 
    12'h970 : errs =          63'b000000000000000000000010000000000000000000100000000000000000000; // D (0x0000010000100000) 
    12'h3d6 : errs =          63'b000000000000000000000010000000000000000001000000000000000000000; // D (0x0000010000200000) 
    12'h3a3 : errs =          63'b000000000000000000000010000000000000000010000000000000000000000; // D (0x0000010000400000) 
    12'h349 : errs =          63'b000000000000000000000010000000000000000100000000000000000000000; // D (0x0000010000800000) 
    12'h29d : errs =          63'b000000000000000000000010000000000000001000000000000000000000000; // D (0x0000010001000000) 
    12'h135 : errs =          63'b000000000000000000000010000000000000010000000000000000000000000; // D (0x0000010002000000) 
    12'h665 : errs =          63'b000000000000000000000010000000000000100000000000000000000000000; // D (0x0000010004000000) 
    12'h8c5 : errs =          63'b000000000000000000000010000000000001000000000000000000000000000; // D (0x0000010008000000) 
    12'h0bc : errs =          63'b000000000000000000000010000000000010000000000000000000000000000; // D (0x0000010010000000) 
    12'h577 : errs =          63'b000000000000000000000010000000000100000000000000000000000000000; // D (0x0000010020000000) 
    12'hee1 : errs =          63'b000000000000000000000010000000001000000000000000000000000000000; // D (0x0000010040000000) 
    12'hcf4 : errs =          63'b000000000000000000000010000000010000000000000000000000000000000; // D (0x0000010080000000) 
    12'h8de : errs =          63'b000000000000000000000010000000100000000000000000000000000000000; // D (0x0000010100000000) 
    12'h08a : errs =          63'b000000000000000000000010000001000000000000000000000000000000000; // D (0x0000010200000000) 
    12'h51b : errs =          63'b000000000000000000000010000010000000000000000000000000000000000; // D (0x0000010400000000) 
    12'he39 : errs =          63'b000000000000000000000010000100000000000000000000000000000000000; // D (0x0000010800000000) 
    12'hd44 : errs =          63'b000000000000000000000010001000000000000000000000000000000000000; // D (0x0000011000000000) 
    12'hbbe : errs =          63'b000000000000000000000010010000000000000000000000000000000000000; // D (0x0000012000000000) 
    12'h64a : errs =          63'b000000000000000000000010100000000000000000000000000000000000000; // D (0x0000014000000000) 
    12'h89b : errs =          63'b000000000000000000000011000000000000000000000000000000000000000; // D (0x0000018000000000) 
    12'hf12 : errs =          63'b000000000000000000000010000000000000000000000000000000000000000; // S (0x0000010000000000) 
//    12'h40f : errs =          63'b000000000000000000000110000000000000000000000000000000000000000; // D (0x0000030000000000) 
//    12'hc11 : errs =          63'b000000000000000000001010000000000000000000000000000000000000000; // D (0x0000050000000000) 
//    12'h914 : errs =          63'b000000000000000000010010000000000000000000000000000000000000000; // D (0x0000090000000000) 
//    12'h31e : errs =          63'b000000000000000000100010000000000000000000000000000000000000000; // D (0x0000110000000000) 
//    12'h233 : errs =          63'b000000000000000001000010000000000000000000000000000000000000000; // D (0x0000210000000000) 
//    12'h069 : errs =          63'b000000000000000010000010000000000000000000000000000000000000000; // D (0x0000410000000000) 
//    12'h4dd : errs =          63'b000000000000000100000010000000000000000000000000000000000000000; // D (0x0000810000000000) 
//    12'hdb5 : errs =          63'b000000000000001000000010000000000000000000000000000000000000000; // D (0x0001010000000000) 
//    12'ha5c : errs =          63'b000000000000010000000010000000000000000000000000000000000000000; // D (0x0002010000000000) 
//    12'h58e : errs =          63'b000000000000100000000010000000000000000000000000000000000000000; // D (0x0004010000000000) 
//    12'hf13 : errs =          63'b000000000001000000000010000000000000000000000000000000000000000; // D (0x0008010000000000) 
//    12'hf10 : errs =          63'b000000000010000000000010000000000000000000000000000000000000000; // D (0x0010010000000000) 
//    12'hf16 : errs =          63'b000000000100000000000010000000000000000000000000000000000000000; // D (0x0020010000000000) 
//    12'hf1a : errs =          63'b000000001000000000000010000000000000000000000000000000000000000; // D (0x0040010000000000) 
//    12'hf02 : errs =          63'b000000010000000000000010000000000000000000000000000000000000000; // D (0x0080010000000000) 
//    12'hf32 : errs =          63'b000000100000000000000010000000000000000000000000000000000000000; // D (0x0100010000000000) 
//    12'hf52 : errs =          63'b000001000000000000000010000000000000000000000000000000000000000; // D (0x0200010000000000) 
//    12'hf92 : errs =          63'b000010000000000000000010000000000000000000000000000000000000000; // D (0x0400010000000000) 
//    12'he12 : errs =          63'b000100000000000000000010000000000000000000000000000000000000000; // D (0x0800010000000000) 
//    12'hd12 : errs =          63'b001000000000000000000010000000000000000000000000000000000000000; // D (0x1000010000000000) 
//    12'hb12 : errs =          63'b010000000000000000000010000000000000000000000000000000000000000; // D (0x2000010000000000) 
//    12'h712 : errs =          63'b100000000000000000000010000000000000000000000000000000000000000; // D (0x4000010000000000) 
    12'he24 : errs =          63'b000000000000000000000100000000000000000000000000000000000000001; // D (0x0000020000000001) 
    12'h16f : errs =          63'b000000000000000000000100000000000000000000000000000000000000010; // D (0x0000020000000002) 
    12'hac0 : errs =          63'b000000000000000000000100000000000000000000000000000000000000100; // D (0x0000020000000004) 
    12'h8a7 : errs =          63'b000000000000000000000100000000000000000000000000000000000001000; // D (0x0000020000000008) 
    12'hc69 : errs =          63'b000000000000000000000100000000000000000000000000000000000010000; // D (0x0000020000000010) 
    12'h5f5 : errs =          63'b000000000000000000000100000000000000000000000000000000000100000; // D (0x0000020000000020) 
    12'h3f4 : errs =          63'b000000000000000000000100000000000000000000000000000000001000000; // D (0x0000020000000040) 
    12'hff6 : errs =          63'b000000000000000000000100000000000000000000000000000000010000000; // D (0x0000020000000080) 
    12'h2cb : errs =          63'b000000000000000000000100000000000000000000000000000000100000000; // D (0x0000020000000100) 
    12'hd88 : errs =          63'b000000000000000000000100000000000000000000000000000001000000000; // D (0x0000020000000200) 
    12'h637 : errs =          63'b000000000000000000000100000000000000000000000000000010000000000; // D (0x0000020000000400) 
    12'h470 : errs =          63'b000000000000000000000100000000000000000000000000000100000000000; // D (0x0000020000000800) 
    12'h0fe : errs =          63'b000000000000000000000100000000000000000000000000001000000000000; // D (0x0000020000001000) 
    12'h9e2 : errs =          63'b000000000000000000000100000000000000000000000000010000000000000; // D (0x0000020000002000) 
    12'hee3 : errs =          63'b000000000000000000000100000000000000000000000000100000000000000; // D (0x0000020000004000) 
    12'h0e1 : errs =          63'b000000000000000000000100000000000000000000000001000000000000000; // D (0x0000020000008000) 
    12'h9dc : errs =          63'b000000000000000000000100000000000000000000000010000000000000000; // D (0x0000020000010000) 
    12'he9f : errs =          63'b000000000000000000000100000000000000000000000100000000000000000; // D (0x0000020000020000) 
    12'h019 : errs =          63'b000000000000000000000100000000000000000000001000000000000000000; // D (0x0000020000040000) 
    12'h82c : errs =          63'b000000000000000000000100000000000000000000010000000000000000000; // D (0x0000020000080000) 
    12'hd7f : errs =          63'b000000000000000000000100000000000000000000100000000000000000000; // D (0x0000020000100000) 
    12'h7d9 : errs =          63'b000000000000000000000100000000000000000001000000000000000000000; // D (0x0000020000200000) 
    12'h7ac : errs =          63'b000000000000000000000100000000000000000010000000000000000000000; // D (0x0000020000400000) 
    12'h746 : errs =          63'b000000000000000000000100000000000000000100000000000000000000000; // D (0x0000020000800000) 
    12'h692 : errs =          63'b000000000000000000000100000000000000001000000000000000000000000; // D (0x0000020001000000) 
    12'h53a : errs =          63'b000000000000000000000100000000000000010000000000000000000000000; // D (0x0000020002000000) 
    12'h26a : errs =          63'b000000000000000000000100000000000000100000000000000000000000000; // D (0x0000020004000000) 
    12'hcca : errs =          63'b000000000000000000000100000000000001000000000000000000000000000; // D (0x0000020008000000) 
    12'h4b3 : errs =          63'b000000000000000000000100000000000010000000000000000000000000000; // D (0x0000020010000000) 
    12'h178 : errs =          63'b000000000000000000000100000000000100000000000000000000000000000; // D (0x0000020020000000) 
    12'haee : errs =          63'b000000000000000000000100000000001000000000000000000000000000000; // D (0x0000020040000000) 
    12'h8fb : errs =          63'b000000000000000000000100000000010000000000000000000000000000000; // D (0x0000020080000000) 
    12'hcd1 : errs =          63'b000000000000000000000100000000100000000000000000000000000000000; // D (0x0000020100000000) 
    12'h485 : errs =          63'b000000000000000000000100000001000000000000000000000000000000000; // D (0x0000020200000000) 
    12'h114 : errs =          63'b000000000000000000000100000010000000000000000000000000000000000; // D (0x0000020400000000) 
    12'ha36 : errs =          63'b000000000000000000000100000100000000000000000000000000000000000; // D (0x0000020800000000) 
    12'h94b : errs =          63'b000000000000000000000100001000000000000000000000000000000000000; // D (0x0000021000000000) 
    12'hfb1 : errs =          63'b000000000000000000000100010000000000000000000000000000000000000; // D (0x0000022000000000) 
    12'h245 : errs =          63'b000000000000000000000100100000000000000000000000000000000000000; // D (0x0000024000000000) 
    12'hc94 : errs =          63'b000000000000000000000101000000000000000000000000000000000000000; // D (0x0000028000000000) 
    12'h40f : errs =          63'b000000000000000000000110000000000000000000000000000000000000000; // D (0x0000030000000000) 
    12'hb1d : errs =          63'b000000000000000000000100000000000000000000000000000000000000000; // S (0x0000020000000000) 
//    12'h81e : errs =          63'b000000000000000000001100000000000000000000000000000000000000000; // D (0x0000060000000000) 
//    12'hd1b : errs =          63'b000000000000000000010100000000000000000000000000000000000000000; // D (0x00000a0000000000) 
//    12'h711 : errs =          63'b000000000000000000100100000000000000000000000000000000000000000; // D (0x0000120000000000) 
//    12'h63c : errs =          63'b000000000000000001000100000000000000000000000000000000000000000; // D (0x0000220000000000) 
//    12'h466 : errs =          63'b000000000000000010000100000000000000000000000000000000000000000; // D (0x0000420000000000) 
//    12'h0d2 : errs =          63'b000000000000000100000100000000000000000000000000000000000000000; // D (0x0000820000000000) 
//    12'h9ba : errs =          63'b000000000000001000000100000000000000000000000000000000000000000; // D (0x0001020000000000) 
//    12'he53 : errs =          63'b000000000000010000000100000000000000000000000000000000000000000; // D (0x0002020000000000) 
//    12'h181 : errs =          63'b000000000000100000000100000000000000000000000000000000000000000; // D (0x0004020000000000) 
//    12'hb1c : errs =          63'b000000000001000000000100000000000000000000000000000000000000000; // D (0x0008020000000000) 
//    12'hb1f : errs =          63'b000000000010000000000100000000000000000000000000000000000000000; // D (0x0010020000000000) 
//    12'hb19 : errs =          63'b000000000100000000000100000000000000000000000000000000000000000; // D (0x0020020000000000) 
//    12'hb15 : errs =          63'b000000001000000000000100000000000000000000000000000000000000000; // D (0x0040020000000000) 
//    12'hb0d : errs =          63'b000000010000000000000100000000000000000000000000000000000000000; // D (0x0080020000000000) 
//    12'hb3d : errs =          63'b000000100000000000000100000000000000000000000000000000000000000; // D (0x0100020000000000) 
//    12'hb5d : errs =          63'b000001000000000000000100000000000000000000000000000000000000000; // D (0x0200020000000000) 
//    12'hb9d : errs =          63'b000010000000000000000100000000000000000000000000000000000000000; // D (0x0400020000000000) 
//    12'ha1d : errs =          63'b000100000000000000000100000000000000000000000000000000000000000; // D (0x0800020000000000) 
//    12'h91d : errs =          63'b001000000000000000000100000000000000000000000000000000000000000; // D (0x1000020000000000) 
//    12'hf1d : errs =          63'b010000000000000000000100000000000000000000000000000000000000000; // D (0x2000020000000000) 
//    12'h31d : errs =          63'b100000000000000000000100000000000000000000000000000000000000000; // D (0x4000020000000000) 
    12'h63a : errs =          63'b000000000000000000001000000000000000000000000000000000000000001; // D (0x0000040000000001) 
    12'h971 : errs =          63'b000000000000000000001000000000000000000000000000000000000000010; // D (0x0000040000000002) 
    12'h2de : errs =          63'b000000000000000000001000000000000000000000000000000000000000100; // D (0x0000040000000004) 
    12'h0b9 : errs =          63'b000000000000000000001000000000000000000000000000000000000001000; // D (0x0000040000000008) 
    12'h477 : errs =          63'b000000000000000000001000000000000000000000000000000000000010000; // D (0x0000040000000010) 
    12'hdeb : errs =          63'b000000000000000000001000000000000000000000000000000000000100000; // D (0x0000040000000020) 
    12'hbea : errs =          63'b000000000000000000001000000000000000000000000000000000001000000; // D (0x0000040000000040) 
    12'h7e8 : errs =          63'b000000000000000000001000000000000000000000000000000000010000000; // D (0x0000040000000080) 
    12'had5 : errs =          63'b000000000000000000001000000000000000000000000000000000100000000; // D (0x0000040000000100) 
    12'h596 : errs =          63'b000000000000000000001000000000000000000000000000000001000000000; // D (0x0000040000000200) 
    12'he29 : errs =          63'b000000000000000000001000000000000000000000000000000010000000000; // D (0x0000040000000400) 
    12'hc6e : errs =          63'b000000000000000000001000000000000000000000000000000100000000000; // D (0x0000040000000800) 
    12'h8e0 : errs =          63'b000000000000000000001000000000000000000000000000001000000000000; // D (0x0000040000001000) 
    12'h1fc : errs =          63'b000000000000000000001000000000000000000000000000010000000000000; // D (0x0000040000002000) 
    12'h6fd : errs =          63'b000000000000000000001000000000000000000000000000100000000000000; // D (0x0000040000004000) 
    12'h8ff : errs =          63'b000000000000000000001000000000000000000000000001000000000000000; // D (0x0000040000008000) 
    12'h1c2 : errs =          63'b000000000000000000001000000000000000000000000010000000000000000; // D (0x0000040000010000) 
    12'h681 : errs =          63'b000000000000000000001000000000000000000000000100000000000000000; // D (0x0000040000020000) 
    12'h807 : errs =          63'b000000000000000000001000000000000000000000001000000000000000000; // D (0x0000040000040000) 
    12'h032 : errs =          63'b000000000000000000001000000000000000000000010000000000000000000; // D (0x0000040000080000) 
    12'h561 : errs =          63'b000000000000000000001000000000000000000000100000000000000000000; // D (0x0000040000100000) 
    12'hfc7 : errs =          63'b000000000000000000001000000000000000000001000000000000000000000; // D (0x0000040000200000) 
    12'hfb2 : errs =          63'b000000000000000000001000000000000000000010000000000000000000000; // D (0x0000040000400000) 
    12'hf58 : errs =          63'b000000000000000000001000000000000000000100000000000000000000000; // D (0x0000040000800000) 
    12'he8c : errs =          63'b000000000000000000001000000000000000001000000000000000000000000; // D (0x0000040001000000) 
    12'hd24 : errs =          63'b000000000000000000001000000000000000010000000000000000000000000; // D (0x0000040002000000) 
    12'ha74 : errs =          63'b000000000000000000001000000000000000100000000000000000000000000; // D (0x0000040004000000) 
    12'h4d4 : errs =          63'b000000000000000000001000000000000001000000000000000000000000000; // D (0x0000040008000000) 
    12'hcad : errs =          63'b000000000000000000001000000000000010000000000000000000000000000; // D (0x0000040010000000) 
    12'h966 : errs =          63'b000000000000000000001000000000000100000000000000000000000000000; // D (0x0000040020000000) 
    12'h2f0 : errs =          63'b000000000000000000001000000000001000000000000000000000000000000; // D (0x0000040040000000) 
    12'h0e5 : errs =          63'b000000000000000000001000000000010000000000000000000000000000000; // D (0x0000040080000000) 
    12'h4cf : errs =          63'b000000000000000000001000000000100000000000000000000000000000000; // D (0x0000040100000000) 
    12'hc9b : errs =          63'b000000000000000000001000000001000000000000000000000000000000000; // D (0x0000040200000000) 
    12'h90a : errs =          63'b000000000000000000001000000010000000000000000000000000000000000; // D (0x0000040400000000) 
    12'h228 : errs =          63'b000000000000000000001000000100000000000000000000000000000000000; // D (0x0000040800000000) 
    12'h155 : errs =          63'b000000000000000000001000001000000000000000000000000000000000000; // D (0x0000041000000000) 
    12'h7af : errs =          63'b000000000000000000001000010000000000000000000000000000000000000; // D (0x0000042000000000) 
    12'ha5b : errs =          63'b000000000000000000001000100000000000000000000000000000000000000; // D (0x0000044000000000) 
    12'h48a : errs =          63'b000000000000000000001001000000000000000000000000000000000000000; // D (0x0000048000000000) 
    12'hc11 : errs =          63'b000000000000000000001010000000000000000000000000000000000000000; // D (0x0000050000000000) 
    12'h81e : errs =          63'b000000000000000000001100000000000000000000000000000000000000000; // D (0x0000060000000000) 
    12'h303 : errs =          63'b000000000000000000001000000000000000000000000000000000000000000; // S (0x0000040000000000) 
//    12'h505 : errs =          63'b000000000000000000011000000000000000000000000000000000000000000; // D (0x00000c0000000000) 
//    12'hf0f : errs =          63'b000000000000000000101000000000000000000000000000000000000000000; // D (0x0000140000000000) 
//    12'he22 : errs =          63'b000000000000000001001000000000000000000000000000000000000000000; // D (0x0000240000000000) 
//    12'hc78 : errs =          63'b000000000000000010001000000000000000000000000000000000000000000; // D (0x0000440000000000) 
//    12'h8cc : errs =          63'b000000000000000100001000000000000000000000000000000000000000000; // D (0x0000840000000000) 
//    12'h1a4 : errs =          63'b000000000000001000001000000000000000000000000000000000000000000; // D (0x0001040000000000) 
//    12'h64d : errs =          63'b000000000000010000001000000000000000000000000000000000000000000; // D (0x0002040000000000) 
//    12'h99f : errs =          63'b000000000000100000001000000000000000000000000000000000000000000; // D (0x0004040000000000) 
//    12'h302 : errs =          63'b000000000001000000001000000000000000000000000000000000000000000; // D (0x0008040000000000) 
//    12'h301 : errs =          63'b000000000010000000001000000000000000000000000000000000000000000; // D (0x0010040000000000) 
//    12'h307 : errs =          63'b000000000100000000001000000000000000000000000000000000000000000; // D (0x0020040000000000) 
//    12'h30b : errs =          63'b000000001000000000001000000000000000000000000000000000000000000; // D (0x0040040000000000) 
//    12'h313 : errs =          63'b000000010000000000001000000000000000000000000000000000000000000; // D (0x0080040000000000) 
//    12'h323 : errs =          63'b000000100000000000001000000000000000000000000000000000000000000; // D (0x0100040000000000) 
//    12'h343 : errs =          63'b000001000000000000001000000000000000000000000000000000000000000; // D (0x0200040000000000) 
//    12'h383 : errs =          63'b000010000000000000001000000000000000000000000000000000000000000; // D (0x0400040000000000) 
//    12'h203 : errs =          63'b000100000000000000001000000000000000000000000000000000000000000; // D (0x0800040000000000) 
//    12'h103 : errs =          63'b001000000000000000001000000000000000000000000000000000000000000; // D (0x1000040000000000) 
//    12'h703 : errs =          63'b010000000000000000001000000000000000000000000000000000000000000; // D (0x2000040000000000) 
//    12'hb03 : errs =          63'b100000000000000000001000000000000000000000000000000000000000000; // D (0x4000040000000000) 
    12'h33f : errs =          63'b000000000000000000010000000000000000000000000000000000000000001; // D (0x0000080000000001) 
    12'hc74 : errs =          63'b000000000000000000010000000000000000000000000000000000000000010; // D (0x0000080000000002) 
    12'h7db : errs =          63'b000000000000000000010000000000000000000000000000000000000000100; // D (0x0000080000000004) 
    12'h5bc : errs =          63'b000000000000000000010000000000000000000000000000000000000001000; // D (0x0000080000000008) 
    12'h172 : errs =          63'b000000000000000000010000000000000000000000000000000000000010000; // D (0x0000080000000010) 
    12'h8ee : errs =          63'b000000000000000000010000000000000000000000000000000000000100000; // D (0x0000080000000020) 
    12'heef : errs =          63'b000000000000000000010000000000000000000000000000000000001000000; // D (0x0000080000000040) 
    12'h2ed : errs =          63'b000000000000000000010000000000000000000000000000000000010000000; // D (0x0000080000000080) 
    12'hfd0 : errs =          63'b000000000000000000010000000000000000000000000000000000100000000; // D (0x0000080000000100) 
    12'h093 : errs =          63'b000000000000000000010000000000000000000000000000000001000000000; // D (0x0000080000000200) 
    12'hb2c : errs =          63'b000000000000000000010000000000000000000000000000000010000000000; // D (0x0000080000000400) 
    12'h96b : errs =          63'b000000000000000000010000000000000000000000000000000100000000000; // D (0x0000080000000800) 
    12'hde5 : errs =          63'b000000000000000000010000000000000000000000000000001000000000000; // D (0x0000080000001000) 
    12'h4f9 : errs =          63'b000000000000000000010000000000000000000000000000010000000000000; // D (0x0000080000002000) 
    12'h3f8 : errs =          63'b000000000000000000010000000000000000000000000000100000000000000; // D (0x0000080000004000) 
    12'hdfa : errs =          63'b000000000000000000010000000000000000000000000001000000000000000; // D (0x0000080000008000) 
    12'h4c7 : errs =          63'b000000000000000000010000000000000000000000000010000000000000000; // D (0x0000080000010000) 
    12'h384 : errs =          63'b000000000000000000010000000000000000000000000100000000000000000; // D (0x0000080000020000) 
    12'hd02 : errs =          63'b000000000000000000010000000000000000000000001000000000000000000; // D (0x0000080000040000) 
    12'h537 : errs =          63'b000000000000000000010000000000000000000000010000000000000000000; // D (0x0000080000080000) 
    12'h064 : errs =          63'b000000000000000000010000000000000000000000100000000000000000000; // D (0x0000080000100000) 
    12'hac2 : errs =          63'b000000000000000000010000000000000000000001000000000000000000000; // D (0x0000080000200000) 
    12'hab7 : errs =          63'b000000000000000000010000000000000000000010000000000000000000000; // D (0x0000080000400000) 
    12'ha5d : errs =          63'b000000000000000000010000000000000000000100000000000000000000000; // D (0x0000080000800000) 
    12'hb89 : errs =          63'b000000000000000000010000000000000000001000000000000000000000000; // D (0x0000080001000000) 
    12'h821 : errs =          63'b000000000000000000010000000000000000010000000000000000000000000; // D (0x0000080002000000) 
    12'hf71 : errs =          63'b000000000000000000010000000000000000100000000000000000000000000; // D (0x0000080004000000) 
    12'h1d1 : errs =          63'b000000000000000000010000000000000001000000000000000000000000000; // D (0x0000080008000000) 
    12'h9a8 : errs =          63'b000000000000000000010000000000000010000000000000000000000000000; // D (0x0000080010000000) 
    12'hc63 : errs =          63'b000000000000000000010000000000000100000000000000000000000000000; // D (0x0000080020000000) 
    12'h7f5 : errs =          63'b000000000000000000010000000000001000000000000000000000000000000; // D (0x0000080040000000) 
    12'h5e0 : errs =          63'b000000000000000000010000000000010000000000000000000000000000000; // D (0x0000080080000000) 
    12'h1ca : errs =          63'b000000000000000000010000000000100000000000000000000000000000000; // D (0x0000080100000000) 
    12'h99e : errs =          63'b000000000000000000010000000001000000000000000000000000000000000; // D (0x0000080200000000) 
    12'hc0f : errs =          63'b000000000000000000010000000010000000000000000000000000000000000; // D (0x0000080400000000) 
    12'h72d : errs =          63'b000000000000000000010000000100000000000000000000000000000000000; // D (0x0000080800000000) 
    12'h450 : errs =          63'b000000000000000000010000001000000000000000000000000000000000000; // D (0x0000081000000000) 
    12'h2aa : errs =          63'b000000000000000000010000010000000000000000000000000000000000000; // D (0x0000082000000000) 
    12'hf5e : errs =          63'b000000000000000000010000100000000000000000000000000000000000000; // D (0x0000084000000000) 
    12'h18f : errs =          63'b000000000000000000010001000000000000000000000000000000000000000; // D (0x0000088000000000) 
    12'h914 : errs =          63'b000000000000000000010010000000000000000000000000000000000000000; // D (0x0000090000000000) 
    12'hd1b : errs =          63'b000000000000000000010100000000000000000000000000000000000000000; // D (0x00000a0000000000) 
    12'h505 : errs =          63'b000000000000000000011000000000000000000000000000000000000000000; // D (0x00000c0000000000) 
    12'h606 : errs =          63'b000000000000000000010000000000000000000000000000000000000000000; // S (0x0000080000000000) 
//    12'ha0a : errs =          63'b000000000000000000110000000000000000000000000000000000000000000; // D (0x0000180000000000) 
//    12'hb27 : errs =          63'b000000000000000001010000000000000000000000000000000000000000000; // D (0x0000280000000000) 
//    12'h97d : errs =          63'b000000000000000010010000000000000000000000000000000000000000000; // D (0x0000480000000000) 
//    12'hdc9 : errs =          63'b000000000000000100010000000000000000000000000000000000000000000; // D (0x0000880000000000) 
//    12'h4a1 : errs =          63'b000000000000001000010000000000000000000000000000000000000000000; // D (0x0001080000000000) 
//    12'h348 : errs =          63'b000000000000010000010000000000000000000000000000000000000000000; // D (0x0002080000000000) 
//    12'hc9a : errs =          63'b000000000000100000010000000000000000000000000000000000000000000; // D (0x0004080000000000) 
//    12'h607 : errs =          63'b000000000001000000010000000000000000000000000000000000000000000; // D (0x0008080000000000) 
//    12'h604 : errs =          63'b000000000010000000010000000000000000000000000000000000000000000; // D (0x0010080000000000) 
//    12'h602 : errs =          63'b000000000100000000010000000000000000000000000000000000000000000; // D (0x0020080000000000) 
//    12'h60e : errs =          63'b000000001000000000010000000000000000000000000000000000000000000; // D (0x0040080000000000) 
//    12'h616 : errs =          63'b000000010000000000010000000000000000000000000000000000000000000; // D (0x0080080000000000) 
//    12'h626 : errs =          63'b000000100000000000010000000000000000000000000000000000000000000; // D (0x0100080000000000) 
//    12'h646 : errs =          63'b000001000000000000010000000000000000000000000000000000000000000; // D (0x0200080000000000) 
//    12'h686 : errs =          63'b000010000000000000010000000000000000000000000000000000000000000; // D (0x0400080000000000) 
//    12'h706 : errs =          63'b000100000000000000010000000000000000000000000000000000000000000; // D (0x0800080000000000) 
//    12'h406 : errs =          63'b001000000000000000010000000000000000000000000000000000000000000; // D (0x1000080000000000) 
//    12'h206 : errs =          63'b010000000000000000010000000000000000000000000000000000000000000; // D (0x2000080000000000) 
//    12'he06 : errs =          63'b100000000000000000010000000000000000000000000000000000000000000; // D (0x4000080000000000) 
    12'h935 : errs =          63'b000000000000000000100000000000000000000000000000000000000000001; // D (0x0000100000000001) 
    12'h67e : errs =          63'b000000000000000000100000000000000000000000000000000000000000010; // D (0x0000100000000002) 
    12'hdd1 : errs =          63'b000000000000000000100000000000000000000000000000000000000000100; // D (0x0000100000000004) 
    12'hfb6 : errs =          63'b000000000000000000100000000000000000000000000000000000000001000; // D (0x0000100000000008) 
    12'hb78 : errs =          63'b000000000000000000100000000000000000000000000000000000000010000; // D (0x0000100000000010) 
    12'h2e4 : errs =          63'b000000000000000000100000000000000000000000000000000000000100000; // D (0x0000100000000020) 
    12'h4e5 : errs =          63'b000000000000000000100000000000000000000000000000000000001000000; // D (0x0000100000000040) 
    12'h8e7 : errs =          63'b000000000000000000100000000000000000000000000000000000010000000; // D (0x0000100000000080) 
    12'h5da : errs =          63'b000000000000000000100000000000000000000000000000000000100000000; // D (0x0000100000000100) 
    12'ha99 : errs =          63'b000000000000000000100000000000000000000000000000000001000000000; // D (0x0000100000000200) 
    12'h126 : errs =          63'b000000000000000000100000000000000000000000000000000010000000000; // D (0x0000100000000400) 
    12'h361 : errs =          63'b000000000000000000100000000000000000000000000000000100000000000; // D (0x0000100000000800) 
    12'h7ef : errs =          63'b000000000000000000100000000000000000000000000000001000000000000; // D (0x0000100000001000) 
    12'hef3 : errs =          63'b000000000000000000100000000000000000000000000000010000000000000; // D (0x0000100000002000) 
    12'h9f2 : errs =          63'b000000000000000000100000000000000000000000000000100000000000000; // D (0x0000100000004000) 
    12'h7f0 : errs =          63'b000000000000000000100000000000000000000000000001000000000000000; // D (0x0000100000008000) 
    12'hecd : errs =          63'b000000000000000000100000000000000000000000000010000000000000000; // D (0x0000100000010000) 
    12'h98e : errs =          63'b000000000000000000100000000000000000000000000100000000000000000; // D (0x0000100000020000) 
    12'h708 : errs =          63'b000000000000000000100000000000000000000000001000000000000000000; // D (0x0000100000040000) 
    12'hf3d : errs =          63'b000000000000000000100000000000000000000000010000000000000000000; // D (0x0000100000080000) 
    12'ha6e : errs =          63'b000000000000000000100000000000000000000000100000000000000000000; // D (0x0000100000100000) 
    12'h0c8 : errs =          63'b000000000000000000100000000000000000000001000000000000000000000; // D (0x0000100000200000) 
    12'h0bd : errs =          63'b000000000000000000100000000000000000000010000000000000000000000; // D (0x0000100000400000) 
    12'h057 : errs =          63'b000000000000000000100000000000000000000100000000000000000000000; // D (0x0000100000800000) 
    12'h183 : errs =          63'b000000000000000000100000000000000000001000000000000000000000000; // D (0x0000100001000000) 
    12'h22b : errs =          63'b000000000000000000100000000000000000010000000000000000000000000; // D (0x0000100002000000) 
    12'h57b : errs =          63'b000000000000000000100000000000000000100000000000000000000000000; // D (0x0000100004000000) 
    12'hbdb : errs =          63'b000000000000000000100000000000000001000000000000000000000000000; // D (0x0000100008000000) 
    12'h3a2 : errs =          63'b000000000000000000100000000000000010000000000000000000000000000; // D (0x0000100010000000) 
    12'h669 : errs =          63'b000000000000000000100000000000000100000000000000000000000000000; // D (0x0000100020000000) 
    12'hdff : errs =          63'b000000000000000000100000000000001000000000000000000000000000000; // D (0x0000100040000000) 
    12'hfea : errs =          63'b000000000000000000100000000000010000000000000000000000000000000; // D (0x0000100080000000) 
    12'hbc0 : errs =          63'b000000000000000000100000000000100000000000000000000000000000000; // D (0x0000100100000000) 
    12'h394 : errs =          63'b000000000000000000100000000001000000000000000000000000000000000; // D (0x0000100200000000) 
    12'h605 : errs =          63'b000000000000000000100000000010000000000000000000000000000000000; // D (0x0000100400000000) 
    12'hd27 : errs =          63'b000000000000000000100000000100000000000000000000000000000000000; // D (0x0000100800000000) 
    12'he5a : errs =          63'b000000000000000000100000001000000000000000000000000000000000000; // D (0x0000101000000000) 
    12'h8a0 : errs =          63'b000000000000000000100000010000000000000000000000000000000000000; // D (0x0000102000000000) 
    12'h554 : errs =          63'b000000000000000000100000100000000000000000000000000000000000000; // D (0x0000104000000000) 
    12'hb85 : errs =          63'b000000000000000000100001000000000000000000000000000000000000000; // D (0x0000108000000000) 
    12'h31e : errs =          63'b000000000000000000100010000000000000000000000000000000000000000; // D (0x0000110000000000) 
    12'h711 : errs =          63'b000000000000000000100100000000000000000000000000000000000000000; // D (0x0000120000000000) 
    12'hf0f : errs =          63'b000000000000000000101000000000000000000000000000000000000000000; // D (0x0000140000000000) 
    12'ha0a : errs =          63'b000000000000000000110000000000000000000000000000000000000000000; // D (0x0000180000000000) 
    12'hc0c : errs =          63'b000000000000000000100000000000000000000000000000000000000000000; // S (0x0000100000000000) 
//    12'h12d : errs =          63'b000000000000000001100000000000000000000000000000000000000000000; // D (0x0000300000000000) 
//    12'h377 : errs =          63'b000000000000000010100000000000000000000000000000000000000000000; // D (0x0000500000000000) 
//    12'h7c3 : errs =          63'b000000000000000100100000000000000000000000000000000000000000000; // D (0x0000900000000000) 
//    12'heab : errs =          63'b000000000000001000100000000000000000000000000000000000000000000; // D (0x0001100000000000) 
//    12'h942 : errs =          63'b000000000000010000100000000000000000000000000000000000000000000; // D (0x0002100000000000) 
//    12'h690 : errs =          63'b000000000000100000100000000000000000000000000000000000000000000; // D (0x0004100000000000) 
//    12'hc0d : errs =          63'b000000000001000000100000000000000000000000000000000000000000000; // D (0x0008100000000000) 
//    12'hc0e : errs =          63'b000000000010000000100000000000000000000000000000000000000000000; // D (0x0010100000000000) 
//    12'hc08 : errs =          63'b000000000100000000100000000000000000000000000000000000000000000; // D (0x0020100000000000) 
//    12'hc04 : errs =          63'b000000001000000000100000000000000000000000000000000000000000000; // D (0x0040100000000000) 
//    12'hc1c : errs =          63'b000000010000000000100000000000000000000000000000000000000000000; // D (0x0080100000000000) 
//    12'hc2c : errs =          63'b000000100000000000100000000000000000000000000000000000000000000; // D (0x0100100000000000) 
//    12'hc4c : errs =          63'b000001000000000000100000000000000000000000000000000000000000000; // D (0x0200100000000000) 
//    12'hc8c : errs =          63'b000010000000000000100000000000000000000000000000000000000000000; // D (0x0400100000000000) 
//    12'hd0c : errs =          63'b000100000000000000100000000000000000000000000000000000000000000; // D (0x0800100000000000) 
//    12'he0c : errs =          63'b001000000000000000100000000000000000000000000000000000000000000; // D (0x1000100000000000) 
//    12'h80c : errs =          63'b010000000000000000100000000000000000000000000000000000000000000; // D (0x2000100000000000) 
//    12'h40c : errs =          63'b100000000000000000100000000000000000000000000000000000000000000; // D (0x4000100000000000) 
    12'h818 : errs =          63'b000000000000000001000000000000000000000000000000000000000000001; // D (0x0000200000000001) 
    12'h753 : errs =          63'b000000000000000001000000000000000000000000000000000000000000010; // D (0x0000200000000002) 
    12'hcfc : errs =          63'b000000000000000001000000000000000000000000000000000000000000100; // D (0x0000200000000004) 
    12'he9b : errs =          63'b000000000000000001000000000000000000000000000000000000000001000; // D (0x0000200000000008) 
    12'ha55 : errs =          63'b000000000000000001000000000000000000000000000000000000000010000; // D (0x0000200000000010) 
    12'h3c9 : errs =          63'b000000000000000001000000000000000000000000000000000000000100000; // D (0x0000200000000020) 
    12'h5c8 : errs =          63'b000000000000000001000000000000000000000000000000000000001000000; // D (0x0000200000000040) 
    12'h9ca : errs =          63'b000000000000000001000000000000000000000000000000000000010000000; // D (0x0000200000000080) 
    12'h4f7 : errs =          63'b000000000000000001000000000000000000000000000000000000100000000; // D (0x0000200000000100) 
    12'hbb4 : errs =          63'b000000000000000001000000000000000000000000000000000001000000000; // D (0x0000200000000200) 
    12'h00b : errs =          63'b000000000000000001000000000000000000000000000000000010000000000; // D (0x0000200000000400) 
    12'h24c : errs =          63'b000000000000000001000000000000000000000000000000000100000000000; // D (0x0000200000000800) 
    12'h6c2 : errs =          63'b000000000000000001000000000000000000000000000000001000000000000; // D (0x0000200000001000) 
    12'hfde : errs =          63'b000000000000000001000000000000000000000000000000010000000000000; // D (0x0000200000002000) 
    12'h8df : errs =          63'b000000000000000001000000000000000000000000000000100000000000000; // D (0x0000200000004000) 
    12'h6dd : errs =          63'b000000000000000001000000000000000000000000000001000000000000000; // D (0x0000200000008000) 
    12'hfe0 : errs =          63'b000000000000000001000000000000000000000000000010000000000000000; // D (0x0000200000010000) 
    12'h8a3 : errs =          63'b000000000000000001000000000000000000000000000100000000000000000; // D (0x0000200000020000) 
    12'h625 : errs =          63'b000000000000000001000000000000000000000000001000000000000000000; // D (0x0000200000040000) 
    12'he10 : errs =          63'b000000000000000001000000000000000000000000010000000000000000000; // D (0x0000200000080000) 
    12'hb43 : errs =          63'b000000000000000001000000000000000000000000100000000000000000000; // D (0x0000200000100000) 
    12'h1e5 : errs =          63'b000000000000000001000000000000000000000001000000000000000000000; // D (0x0000200000200000) 
    12'h190 : errs =          63'b000000000000000001000000000000000000000010000000000000000000000; // D (0x0000200000400000) 
    12'h17a : errs =          63'b000000000000000001000000000000000000000100000000000000000000000; // D (0x0000200000800000) 
    12'h0ae : errs =          63'b000000000000000001000000000000000000001000000000000000000000000; // D (0x0000200001000000) 
    12'h306 : errs =          63'b000000000000000001000000000000000000010000000000000000000000000; // D (0x0000200002000000) 
    12'h456 : errs =          63'b000000000000000001000000000000000000100000000000000000000000000; // D (0x0000200004000000) 
    12'haf6 : errs =          63'b000000000000000001000000000000000001000000000000000000000000000; // D (0x0000200008000000) 
    12'h28f : errs =          63'b000000000000000001000000000000000010000000000000000000000000000; // D (0x0000200010000000) 
    12'h744 : errs =          63'b000000000000000001000000000000000100000000000000000000000000000; // D (0x0000200020000000) 
    12'hcd2 : errs =          63'b000000000000000001000000000000001000000000000000000000000000000; // D (0x0000200040000000) 
    12'hec7 : errs =          63'b000000000000000001000000000000010000000000000000000000000000000; // D (0x0000200080000000) 
    12'haed : errs =          63'b000000000000000001000000000000100000000000000000000000000000000; // D (0x0000200100000000) 
    12'h2b9 : errs =          63'b000000000000000001000000000001000000000000000000000000000000000; // D (0x0000200200000000) 
    12'h728 : errs =          63'b000000000000000001000000000010000000000000000000000000000000000; // D (0x0000200400000000) 
    12'hc0a : errs =          63'b000000000000000001000000000100000000000000000000000000000000000; // D (0x0000200800000000) 
    12'hf77 : errs =          63'b000000000000000001000000001000000000000000000000000000000000000; // D (0x0000201000000000) 
    12'h98d : errs =          63'b000000000000000001000000010000000000000000000000000000000000000; // D (0x0000202000000000) 
    12'h479 : errs =          63'b000000000000000001000000100000000000000000000000000000000000000; // D (0x0000204000000000) 
    12'haa8 : errs =          63'b000000000000000001000001000000000000000000000000000000000000000; // D (0x0000208000000000) 
    12'h233 : errs =          63'b000000000000000001000010000000000000000000000000000000000000000; // D (0x0000210000000000) 
    12'h63c : errs =          63'b000000000000000001000100000000000000000000000000000000000000000; // D (0x0000220000000000) 
    12'he22 : errs =          63'b000000000000000001001000000000000000000000000000000000000000000; // D (0x0000240000000000) 
    12'hb27 : errs =          63'b000000000000000001010000000000000000000000000000000000000000000; // D (0x0000280000000000) 
    12'h12d : errs =          63'b000000000000000001100000000000000000000000000000000000000000000; // D (0x0000300000000000) 
    12'hd21 : errs =          63'b000000000000000001000000000000000000000000000000000000000000000; // S (0x0000200000000000) 
//    12'h25a : errs =          63'b000000000000000011000000000000000000000000000000000000000000000; // D (0x0000600000000000) 
//    12'h6ee : errs =          63'b000000000000000101000000000000000000000000000000000000000000000; // D (0x0000a00000000000) 
//    12'hf86 : errs =          63'b000000000000001001000000000000000000000000000000000000000000000; // D (0x0001200000000000) 
//    12'h86f : errs =          63'b000000000000010001000000000000000000000000000000000000000000000; // D (0x0002200000000000) 
//    12'h7bd : errs =          63'b000000000000100001000000000000000000000000000000000000000000000; // D (0x0004200000000000) 
//    12'hd20 : errs =          63'b000000000001000001000000000000000000000000000000000000000000000; // D (0x0008200000000000) 
//    12'hd23 : errs =          63'b000000000010000001000000000000000000000000000000000000000000000; // D (0x0010200000000000) 
//    12'hd25 : errs =          63'b000000000100000001000000000000000000000000000000000000000000000; // D (0x0020200000000000) 
//    12'hd29 : errs =          63'b000000001000000001000000000000000000000000000000000000000000000; // D (0x0040200000000000) 
//    12'hd31 : errs =          63'b000000010000000001000000000000000000000000000000000000000000000; // D (0x0080200000000000) 
//    12'hd01 : errs =          63'b000000100000000001000000000000000000000000000000000000000000000; // D (0x0100200000000000) 
//    12'hd61 : errs =          63'b000001000000000001000000000000000000000000000000000000000000000; // D (0x0200200000000000) 
//    12'hda1 : errs =          63'b000010000000000001000000000000000000000000000000000000000000000; // D (0x0400200000000000) 
//    12'hc21 : errs =          63'b000100000000000001000000000000000000000000000000000000000000000; // D (0x0800200000000000) 
//    12'hf21 : errs =          63'b001000000000000001000000000000000000000000000000000000000000000; // D (0x1000200000000000) 
//    12'h921 : errs =          63'b010000000000000001000000000000000000000000000000000000000000000; // D (0x2000200000000000) 
//    12'h521 : errs =          63'b100000000000000001000000000000000000000000000000000000000000000; // D (0x4000200000000000) 
    12'ha42 : errs =          63'b000000000000000010000000000000000000000000000000000000000000001; // D (0x0000400000000001) 
    12'h509 : errs =          63'b000000000000000010000000000000000000000000000000000000000000010; // D (0x0000400000000002) 
    12'hea6 : errs =          63'b000000000000000010000000000000000000000000000000000000000000100; // D (0x0000400000000004) 
    12'hcc1 : errs =          63'b000000000000000010000000000000000000000000000000000000000001000; // D (0x0000400000000008) 
    12'h80f : errs =          63'b000000000000000010000000000000000000000000000000000000000010000; // D (0x0000400000000010) 
    12'h193 : errs =          63'b000000000000000010000000000000000000000000000000000000000100000; // D (0x0000400000000020) 
    12'h792 : errs =          63'b000000000000000010000000000000000000000000000000000000001000000; // D (0x0000400000000040) 
    12'hb90 : errs =          63'b000000000000000010000000000000000000000000000000000000010000000; // D (0x0000400000000080) 
    12'h6ad : errs =          63'b000000000000000010000000000000000000000000000000000000100000000; // D (0x0000400000000100) 
    12'h9ee : errs =          63'b000000000000000010000000000000000000000000000000000001000000000; // D (0x0000400000000200) 
    12'h251 : errs =          63'b000000000000000010000000000000000000000000000000000010000000000; // D (0x0000400000000400) 
    12'h016 : errs =          63'b000000000000000010000000000000000000000000000000000100000000000; // D (0x0000400000000800) 
    12'h498 : errs =          63'b000000000000000010000000000000000000000000000000001000000000000; // D (0x0000400000001000) 
    12'hd84 : errs =          63'b000000000000000010000000000000000000000000000000010000000000000; // D (0x0000400000002000) 
    12'ha85 : errs =          63'b000000000000000010000000000000000000000000000000100000000000000; // D (0x0000400000004000) 
    12'h487 : errs =          63'b000000000000000010000000000000000000000000000001000000000000000; // D (0x0000400000008000) 
    12'hdba : errs =          63'b000000000000000010000000000000000000000000000010000000000000000; // D (0x0000400000010000) 
    12'haf9 : errs =          63'b000000000000000010000000000000000000000000000100000000000000000; // D (0x0000400000020000) 
    12'h47f : errs =          63'b000000000000000010000000000000000000000000001000000000000000000; // D (0x0000400000040000) 
    12'hc4a : errs =          63'b000000000000000010000000000000000000000000010000000000000000000; // D (0x0000400000080000) 
    12'h919 : errs =          63'b000000000000000010000000000000000000000000100000000000000000000; // D (0x0000400000100000) 
    12'h3bf : errs =          63'b000000000000000010000000000000000000000001000000000000000000000; // D (0x0000400000200000) 
    12'h3ca : errs =          63'b000000000000000010000000000000000000000010000000000000000000000; // D (0x0000400000400000) 
    12'h320 : errs =          63'b000000000000000010000000000000000000000100000000000000000000000; // D (0x0000400000800000) 
    12'h2f4 : errs =          63'b000000000000000010000000000000000000001000000000000000000000000; // D (0x0000400001000000) 
    12'h15c : errs =          63'b000000000000000010000000000000000000010000000000000000000000000; // D (0x0000400002000000) 
    12'h60c : errs =          63'b000000000000000010000000000000000000100000000000000000000000000; // D (0x0000400004000000) 
    12'h8ac : errs =          63'b000000000000000010000000000000000001000000000000000000000000000; // D (0x0000400008000000) 
    12'h0d5 : errs =          63'b000000000000000010000000000000000010000000000000000000000000000; // D (0x0000400010000000) 
    12'h51e : errs =          63'b000000000000000010000000000000000100000000000000000000000000000; // D (0x0000400020000000) 
    12'he88 : errs =          63'b000000000000000010000000000000001000000000000000000000000000000; // D (0x0000400040000000) 
    12'hc9d : errs =          63'b000000000000000010000000000000010000000000000000000000000000000; // D (0x0000400080000000) 
    12'h8b7 : errs =          63'b000000000000000010000000000000100000000000000000000000000000000; // D (0x0000400100000000) 
    12'h0e3 : errs =          63'b000000000000000010000000000001000000000000000000000000000000000; // D (0x0000400200000000) 
    12'h572 : errs =          63'b000000000000000010000000000010000000000000000000000000000000000; // D (0x0000400400000000) 
    12'he50 : errs =          63'b000000000000000010000000000100000000000000000000000000000000000; // D (0x0000400800000000) 
    12'hd2d : errs =          63'b000000000000000010000000001000000000000000000000000000000000000; // D (0x0000401000000000) 
    12'hbd7 : errs =          63'b000000000000000010000000010000000000000000000000000000000000000; // D (0x0000402000000000) 
    12'h623 : errs =          63'b000000000000000010000000100000000000000000000000000000000000000; // D (0x0000404000000000) 
    12'h8f2 : errs =          63'b000000000000000010000001000000000000000000000000000000000000000; // D (0x0000408000000000) 
    12'h069 : errs =          63'b000000000000000010000010000000000000000000000000000000000000000; // D (0x0000410000000000) 
    12'h466 : errs =          63'b000000000000000010000100000000000000000000000000000000000000000; // D (0x0000420000000000) 
    12'hc78 : errs =          63'b000000000000000010001000000000000000000000000000000000000000000; // D (0x0000440000000000) 
    12'h97d : errs =          63'b000000000000000010010000000000000000000000000000000000000000000; // D (0x0000480000000000) 
    12'h377 : errs =          63'b000000000000000010100000000000000000000000000000000000000000000; // D (0x0000500000000000) 
    12'h25a : errs =          63'b000000000000000011000000000000000000000000000000000000000000000; // D (0x0000600000000000) 
    12'hf7b : errs =          63'b000000000000000010000000000000000000000000000000000000000000000; // S (0x0000400000000000) 
//    12'h4b4 : errs =          63'b000000000000000110000000000000000000000000000000000000000000000; // D (0x0000c00000000000) 
//    12'hddc : errs =          63'b000000000000001010000000000000000000000000000000000000000000000; // D (0x0001400000000000) 
//    12'ha35 : errs =          63'b000000000000010010000000000000000000000000000000000000000000000; // D (0x0002400000000000) 
//    12'h5e7 : errs =          63'b000000000000100010000000000000000000000000000000000000000000000; // D (0x0004400000000000) 
//    12'hf7a : errs =          63'b000000000001000010000000000000000000000000000000000000000000000; // D (0x0008400000000000) 
//    12'hf79 : errs =          63'b000000000010000010000000000000000000000000000000000000000000000; // D (0x0010400000000000) 
//    12'hf7f : errs =          63'b000000000100000010000000000000000000000000000000000000000000000; // D (0x0020400000000000) 
//    12'hf73 : errs =          63'b000000001000000010000000000000000000000000000000000000000000000; // D (0x0040400000000000) 
//    12'hf6b : errs =          63'b000000010000000010000000000000000000000000000000000000000000000; // D (0x0080400000000000) 
//    12'hf5b : errs =          63'b000000100000000010000000000000000000000000000000000000000000000; // D (0x0100400000000000) 
//    12'hf3b : errs =          63'b000001000000000010000000000000000000000000000000000000000000000; // D (0x0200400000000000) 
//    12'hffb : errs =          63'b000010000000000010000000000000000000000000000000000000000000000; // D (0x0400400000000000) 
//    12'he7b : errs =          63'b000100000000000010000000000000000000000000000000000000000000000; // D (0x0800400000000000) 
//    12'hd7b : errs =          63'b001000000000000010000000000000000000000000000000000000000000000; // D (0x1000400000000000) 
//    12'hb7b : errs =          63'b010000000000000010000000000000000000000000000000000000000000000; // D (0x2000400000000000) 
//    12'h77b : errs =          63'b100000000000000010000000000000000000000000000000000000000000000; // D (0x4000400000000000) 
    12'hef6 : errs =          63'b000000000000000100000000000000000000000000000000000000000000001; // D (0x0000800000000001) 
    12'h1bd : errs =          63'b000000000000000100000000000000000000000000000000000000000000010; // D (0x0000800000000002) 
    12'ha12 : errs =          63'b000000000000000100000000000000000000000000000000000000000000100; // D (0x0000800000000004) 
    12'h875 : errs =          63'b000000000000000100000000000000000000000000000000000000000001000; // D (0x0000800000000008) 
    12'hcbb : errs =          63'b000000000000000100000000000000000000000000000000000000000010000; // D (0x0000800000000010) 
    12'h527 : errs =          63'b000000000000000100000000000000000000000000000000000000000100000; // D (0x0000800000000020) 
    12'h326 : errs =          63'b000000000000000100000000000000000000000000000000000000001000000; // D (0x0000800000000040) 
    12'hf24 : errs =          63'b000000000000000100000000000000000000000000000000000000010000000; // D (0x0000800000000080) 
    12'h219 : errs =          63'b000000000000000100000000000000000000000000000000000000100000000; // D (0x0000800000000100) 
    12'hd5a : errs =          63'b000000000000000100000000000000000000000000000000000001000000000; // D (0x0000800000000200) 
    12'h6e5 : errs =          63'b000000000000000100000000000000000000000000000000000010000000000; // D (0x0000800000000400) 
    12'h4a2 : errs =          63'b000000000000000100000000000000000000000000000000000100000000000; // D (0x0000800000000800) 
    12'h02c : errs =          63'b000000000000000100000000000000000000000000000000001000000000000; // D (0x0000800000001000) 
    12'h930 : errs =          63'b000000000000000100000000000000000000000000000000010000000000000; // D (0x0000800000002000) 
    12'he31 : errs =          63'b000000000000000100000000000000000000000000000000100000000000000; // D (0x0000800000004000) 
    12'h033 : errs =          63'b000000000000000100000000000000000000000000000001000000000000000; // D (0x0000800000008000) 
    12'h90e : errs =          63'b000000000000000100000000000000000000000000000010000000000000000; // D (0x0000800000010000) 
    12'he4d : errs =          63'b000000000000000100000000000000000000000000000100000000000000000; // D (0x0000800000020000) 
    12'h0cb : errs =          63'b000000000000000100000000000000000000000000001000000000000000000; // D (0x0000800000040000) 
    12'h8fe : errs =          63'b000000000000000100000000000000000000000000010000000000000000000; // D (0x0000800000080000) 
    12'hdad : errs =          63'b000000000000000100000000000000000000000000100000000000000000000; // D (0x0000800000100000) 
    12'h70b : errs =          63'b000000000000000100000000000000000000000001000000000000000000000; // D (0x0000800000200000) 
    12'h77e : errs =          63'b000000000000000100000000000000000000000010000000000000000000000; // D (0x0000800000400000) 
    12'h794 : errs =          63'b000000000000000100000000000000000000000100000000000000000000000; // D (0x0000800000800000) 
    12'h640 : errs =          63'b000000000000000100000000000000000000001000000000000000000000000; // D (0x0000800001000000) 
    12'h5e8 : errs =          63'b000000000000000100000000000000000000010000000000000000000000000; // D (0x0000800002000000) 
    12'h2b8 : errs =          63'b000000000000000100000000000000000000100000000000000000000000000; // D (0x0000800004000000) 
    12'hc18 : errs =          63'b000000000000000100000000000000000001000000000000000000000000000; // D (0x0000800008000000) 
    12'h461 : errs =          63'b000000000000000100000000000000000010000000000000000000000000000; // D (0x0000800010000000) 
    12'h1aa : errs =          63'b000000000000000100000000000000000100000000000000000000000000000; // D (0x0000800020000000) 
    12'ha3c : errs =          63'b000000000000000100000000000000001000000000000000000000000000000; // D (0x0000800040000000) 
    12'h829 : errs =          63'b000000000000000100000000000000010000000000000000000000000000000; // D (0x0000800080000000) 
    12'hc03 : errs =          63'b000000000000000100000000000000100000000000000000000000000000000; // D (0x0000800100000000) 
    12'h457 : errs =          63'b000000000000000100000000000001000000000000000000000000000000000; // D (0x0000800200000000) 
    12'h1c6 : errs =          63'b000000000000000100000000000010000000000000000000000000000000000; // D (0x0000800400000000) 
    12'hae4 : errs =          63'b000000000000000100000000000100000000000000000000000000000000000; // D (0x0000800800000000) 
    12'h999 : errs =          63'b000000000000000100000000001000000000000000000000000000000000000; // D (0x0000801000000000) 
    12'hf63 : errs =          63'b000000000000000100000000010000000000000000000000000000000000000; // D (0x0000802000000000) 
    12'h297 : errs =          63'b000000000000000100000000100000000000000000000000000000000000000; // D (0x0000804000000000) 
    12'hc46 : errs =          63'b000000000000000100000001000000000000000000000000000000000000000; // D (0x0000808000000000) 
    12'h4dd : errs =          63'b000000000000000100000010000000000000000000000000000000000000000; // D (0x0000810000000000) 
    12'h0d2 : errs =          63'b000000000000000100000100000000000000000000000000000000000000000; // D (0x0000820000000000) 
    12'h8cc : errs =          63'b000000000000000100001000000000000000000000000000000000000000000; // D (0x0000840000000000) 
    12'hdc9 : errs =          63'b000000000000000100010000000000000000000000000000000000000000000; // D (0x0000880000000000) 
    12'h7c3 : errs =          63'b000000000000000100100000000000000000000000000000000000000000000; // D (0x0000900000000000) 
    12'h6ee : errs =          63'b000000000000000101000000000000000000000000000000000000000000000; // D (0x0000a00000000000) 
    12'h4b4 : errs =          63'b000000000000000110000000000000000000000000000000000000000000000; // D (0x0000c00000000000) 
    12'hbcf : errs =          63'b000000000000000100000000000000000000000000000000000000000000000; // S (0x0000800000000000) 
//    12'h968 : errs =          63'b000000000000001100000000000000000000000000000000000000000000000; // D (0x0001800000000000) 
//    12'he81 : errs =          63'b000000000000010100000000000000000000000000000000000000000000000; // D (0x0002800000000000) 
//    12'h153 : errs =          63'b000000000000100100000000000000000000000000000000000000000000000; // D (0x0004800000000000) 
//    12'hbce : errs =          63'b000000000001000100000000000000000000000000000000000000000000000; // D (0x0008800000000000) 
//    12'hbcd : errs =          63'b000000000010000100000000000000000000000000000000000000000000000; // D (0x0010800000000000) 
//    12'hbcb : errs =          63'b000000000100000100000000000000000000000000000000000000000000000; // D (0x0020800000000000) 
//    12'hbc7 : errs =          63'b000000001000000100000000000000000000000000000000000000000000000; // D (0x0040800000000000) 
//    12'hbdf : errs =          63'b000000010000000100000000000000000000000000000000000000000000000; // D (0x0080800000000000) 
//    12'hbef : errs =          63'b000000100000000100000000000000000000000000000000000000000000000; // D (0x0100800000000000) 
//    12'hb8f : errs =          63'b000001000000000100000000000000000000000000000000000000000000000; // D (0x0200800000000000) 
//    12'hb4f : errs =          63'b000010000000000100000000000000000000000000000000000000000000000; // D (0x0400800000000000) 
//    12'hacf : errs =          63'b000100000000000100000000000000000000000000000000000000000000000; // D (0x0800800000000000) 
//    12'h9cf : errs =          63'b001000000000000100000000000000000000000000000000000000000000000; // D (0x1000800000000000) 
//    12'hfcf : errs =          63'b010000000000000100000000000000000000000000000000000000000000000; // D (0x2000800000000000) 
//    12'h3cf : errs =          63'b100000000000000100000000000000000000000000000000000000000000000; // D (0x4000800000000000) 
    12'h79e : errs =          63'b000000000000001000000000000000000000000000000000000000000000001; // D (0x0001000000000001) 
    12'h8d5 : errs =          63'b000000000000001000000000000000000000000000000000000000000000010; // D (0x0001000000000002) 
    12'h37a : errs =          63'b000000000000001000000000000000000000000000000000000000000000100; // D (0x0001000000000004) 
    12'h11d : errs =          63'b000000000000001000000000000000000000000000000000000000000001000; // D (0x0001000000000008) 
    12'h5d3 : errs =          63'b000000000000001000000000000000000000000000000000000000000010000; // D (0x0001000000000010) 
    12'hc4f : errs =          63'b000000000000001000000000000000000000000000000000000000000100000; // D (0x0001000000000020) 
    12'ha4e : errs =          63'b000000000000001000000000000000000000000000000000000000001000000; // D (0x0001000000000040) 
    12'h64c : errs =          63'b000000000000001000000000000000000000000000000000000000010000000; // D (0x0001000000000080) 
    12'hb71 : errs =          63'b000000000000001000000000000000000000000000000000000000100000000; // D (0x0001000000000100) 
    12'h432 : errs =          63'b000000000000001000000000000000000000000000000000000001000000000; // D (0x0001000000000200) 
    12'hf8d : errs =          63'b000000000000001000000000000000000000000000000000000010000000000; // D (0x0001000000000400) 
    12'hdca : errs =          63'b000000000000001000000000000000000000000000000000000100000000000; // D (0x0001000000000800) 
    12'h944 : errs =          63'b000000000000001000000000000000000000000000000000001000000000000; // D (0x0001000000001000) 
    12'h058 : errs =          63'b000000000000001000000000000000000000000000000000010000000000000; // D (0x0001000000002000) 
    12'h759 : errs =          63'b000000000000001000000000000000000000000000000000100000000000000; // D (0x0001000000004000) 
    12'h95b : errs =          63'b000000000000001000000000000000000000000000000001000000000000000; // D (0x0001000000008000) 
    12'h066 : errs =          63'b000000000000001000000000000000000000000000000010000000000000000; // D (0x0001000000010000) 
    12'h725 : errs =          63'b000000000000001000000000000000000000000000000100000000000000000; // D (0x0001000000020000) 
    12'h9a3 : errs =          63'b000000000000001000000000000000000000000000001000000000000000000; // D (0x0001000000040000) 
    12'h196 : errs =          63'b000000000000001000000000000000000000000000010000000000000000000; // D (0x0001000000080000) 
    12'h4c5 : errs =          63'b000000000000001000000000000000000000000000100000000000000000000; // D (0x0001000000100000) 
    12'he63 : errs =          63'b000000000000001000000000000000000000000001000000000000000000000; // D (0x0001000000200000) 
    12'he16 : errs =          63'b000000000000001000000000000000000000000010000000000000000000000; // D (0x0001000000400000) 
    12'hefc : errs =          63'b000000000000001000000000000000000000000100000000000000000000000; // D (0x0001000000800000) 
    12'hf28 : errs =          63'b000000000000001000000000000000000000001000000000000000000000000; // D (0x0001000001000000) 
    12'hc80 : errs =          63'b000000000000001000000000000000000000010000000000000000000000000; // D (0x0001000002000000) 
    12'hbd0 : errs =          63'b000000000000001000000000000000000000100000000000000000000000000; // D (0x0001000004000000) 
    12'h570 : errs =          63'b000000000000001000000000000000000001000000000000000000000000000; // D (0x0001000008000000) 
    12'hd09 : errs =          63'b000000000000001000000000000000000010000000000000000000000000000; // D (0x0001000010000000) 
    12'h8c2 : errs =          63'b000000000000001000000000000000000100000000000000000000000000000; // D (0x0001000020000000) 
    12'h354 : errs =          63'b000000000000001000000000000000001000000000000000000000000000000; // D (0x0001000040000000) 
    12'h141 : errs =          63'b000000000000001000000000000000010000000000000000000000000000000; // D (0x0001000080000000) 
    12'h56b : errs =          63'b000000000000001000000000000000100000000000000000000000000000000; // D (0x0001000100000000) 
    12'hd3f : errs =          63'b000000000000001000000000000001000000000000000000000000000000000; // D (0x0001000200000000) 
    12'h8ae : errs =          63'b000000000000001000000000000010000000000000000000000000000000000; // D (0x0001000400000000) 
    12'h38c : errs =          63'b000000000000001000000000000100000000000000000000000000000000000; // D (0x0001000800000000) 
    12'h0f1 : errs =          63'b000000000000001000000000001000000000000000000000000000000000000; // D (0x0001001000000000) 
    12'h60b : errs =          63'b000000000000001000000000010000000000000000000000000000000000000; // D (0x0001002000000000) 
    12'hbff : errs =          63'b000000000000001000000000100000000000000000000000000000000000000; // D (0x0001004000000000) 
    12'h52e : errs =          63'b000000000000001000000001000000000000000000000000000000000000000; // D (0x0001008000000000) 
    12'hdb5 : errs =          63'b000000000000001000000010000000000000000000000000000000000000000; // D (0x0001010000000000) 
    12'h9ba : errs =          63'b000000000000001000000100000000000000000000000000000000000000000; // D (0x0001020000000000) 
    12'h1a4 : errs =          63'b000000000000001000001000000000000000000000000000000000000000000; // D (0x0001040000000000) 
    12'h4a1 : errs =          63'b000000000000001000010000000000000000000000000000000000000000000; // D (0x0001080000000000) 
    12'heab : errs =          63'b000000000000001000100000000000000000000000000000000000000000000; // D (0x0001100000000000) 
    12'hf86 : errs =          63'b000000000000001001000000000000000000000000000000000000000000000; // D (0x0001200000000000) 
    12'hddc : errs =          63'b000000000000001010000000000000000000000000000000000000000000000; // D (0x0001400000000000) 
    12'h968 : errs =          63'b000000000000001100000000000000000000000000000000000000000000000; // D (0x0001800000000000) 
    12'h2a7 : errs =          63'b000000000000001000000000000000000000000000000000000000000000000; // S (0x0001000000000000) 
//    12'h7e9 : errs =          63'b000000000000011000000000000000000000000000000000000000000000000; // D (0x0003000000000000) 
//    12'h83b : errs =          63'b000000000000101000000000000000000000000000000000000000000000000; // D (0x0005000000000000) 
//    12'h2a6 : errs =          63'b000000000001001000000000000000000000000000000000000000000000000; // D (0x0009000000000000) 
//    12'h2a5 : errs =          63'b000000000010001000000000000000000000000000000000000000000000000; // D (0x0011000000000000) 
//    12'h2a3 : errs =          63'b000000000100001000000000000000000000000000000000000000000000000; // D (0x0021000000000000) 
//    12'h2af : errs =          63'b000000001000001000000000000000000000000000000000000000000000000; // D (0x0041000000000000) 
//    12'h2b7 : errs =          63'b000000010000001000000000000000000000000000000000000000000000000; // D (0x0081000000000000) 
//    12'h287 : errs =          63'b000000100000001000000000000000000000000000000000000000000000000; // D (0x0101000000000000) 
//    12'h2e7 : errs =          63'b000001000000001000000000000000000000000000000000000000000000000; // D (0x0201000000000000) 
//    12'h227 : errs =          63'b000010000000001000000000000000000000000000000000000000000000000; // D (0x0401000000000000) 
//    12'h3a7 : errs =          63'b000100000000001000000000000000000000000000000000000000000000000; // D (0x0801000000000000) 
//    12'h0a7 : errs =          63'b001000000000001000000000000000000000000000000000000000000000000; // D (0x1001000000000000) 
//    12'h6a7 : errs =          63'b010000000000001000000000000000000000000000000000000000000000000; // D (0x2001000000000000) 
//    12'haa7 : errs =          63'b100000000000001000000000000000000000000000000000000000000000000; // D (0x4001000000000000) 
    12'h077 : errs =          63'b000000000000010000000000000000000000000000000000000000000000001; // D (0x0002000000000001) 
    12'hf3c : errs =          63'b000000000000010000000000000000000000000000000000000000000000010; // D (0x0002000000000002) 
    12'h493 : errs =          63'b000000000000010000000000000000000000000000000000000000000000100; // D (0x0002000000000004) 
    12'h6f4 : errs =          63'b000000000000010000000000000000000000000000000000000000000001000; // D (0x0002000000000008) 
    12'h23a : errs =          63'b000000000000010000000000000000000000000000000000000000000010000; // D (0x0002000000000010) 
    12'hba6 : errs =          63'b000000000000010000000000000000000000000000000000000000000100000; // D (0x0002000000000020) 
    12'hda7 : errs =          63'b000000000000010000000000000000000000000000000000000000001000000; // D (0x0002000000000040) 
    12'h1a5 : errs =          63'b000000000000010000000000000000000000000000000000000000010000000; // D (0x0002000000000080) 
    12'hc98 : errs =          63'b000000000000010000000000000000000000000000000000000000100000000; // D (0x0002000000000100) 
    12'h3db : errs =          63'b000000000000010000000000000000000000000000000000000001000000000; // D (0x0002000000000200) 
    12'h864 : errs =          63'b000000000000010000000000000000000000000000000000000010000000000; // D (0x0002000000000400) 
    12'ha23 : errs =          63'b000000000000010000000000000000000000000000000000000100000000000; // D (0x0002000000000800) 
    12'head : errs =          63'b000000000000010000000000000000000000000000000000001000000000000; // D (0x0002000000001000) 
    12'h7b1 : errs =          63'b000000000000010000000000000000000000000000000000010000000000000; // D (0x0002000000002000) 
    12'h0b0 : errs =          63'b000000000000010000000000000000000000000000000000100000000000000; // D (0x0002000000004000) 
    12'heb2 : errs =          63'b000000000000010000000000000000000000000000000001000000000000000; // D (0x0002000000008000) 
    12'h78f : errs =          63'b000000000000010000000000000000000000000000000010000000000000000; // D (0x0002000000010000) 
    12'h0cc : errs =          63'b000000000000010000000000000000000000000000000100000000000000000; // D (0x0002000000020000) 
    12'he4a : errs =          63'b000000000000010000000000000000000000000000001000000000000000000; // D (0x0002000000040000) 
    12'h67f : errs =          63'b000000000000010000000000000000000000000000010000000000000000000; // D (0x0002000000080000) 
    12'h32c : errs =          63'b000000000000010000000000000000000000000000100000000000000000000; // D (0x0002000000100000) 
    12'h98a : errs =          63'b000000000000010000000000000000000000000001000000000000000000000; // D (0x0002000000200000) 
    12'h9ff : errs =          63'b000000000000010000000000000000000000000010000000000000000000000; // D (0x0002000000400000) 
    12'h915 : errs =          63'b000000000000010000000000000000000000000100000000000000000000000; // D (0x0002000000800000) 
    12'h8c1 : errs =          63'b000000000000010000000000000000000000001000000000000000000000000; // D (0x0002000001000000) 
    12'hb69 : errs =          63'b000000000000010000000000000000000000010000000000000000000000000; // D (0x0002000002000000) 
    12'hc39 : errs =          63'b000000000000010000000000000000000000100000000000000000000000000; // D (0x0002000004000000) 
    12'h299 : errs =          63'b000000000000010000000000000000000001000000000000000000000000000; // D (0x0002000008000000) 
    12'hae0 : errs =          63'b000000000000010000000000000000000010000000000000000000000000000; // D (0x0002000010000000) 
    12'hf2b : errs =          63'b000000000000010000000000000000000100000000000000000000000000000; // D (0x0002000020000000) 
    12'h4bd : errs =          63'b000000000000010000000000000000001000000000000000000000000000000; // D (0x0002000040000000) 
    12'h6a8 : errs =          63'b000000000000010000000000000000010000000000000000000000000000000; // D (0x0002000080000000) 
    12'h282 : errs =          63'b000000000000010000000000000000100000000000000000000000000000000; // D (0x0002000100000000) 
    12'had6 : errs =          63'b000000000000010000000000000001000000000000000000000000000000000; // D (0x0002000200000000) 
    12'hf47 : errs =          63'b000000000000010000000000000010000000000000000000000000000000000; // D (0x0002000400000000) 
    12'h465 : errs =          63'b000000000000010000000000000100000000000000000000000000000000000; // D (0x0002000800000000) 
    12'h718 : errs =          63'b000000000000010000000000001000000000000000000000000000000000000; // D (0x0002001000000000) 
    12'h1e2 : errs =          63'b000000000000010000000000010000000000000000000000000000000000000; // D (0x0002002000000000) 
    12'hc16 : errs =          63'b000000000000010000000000100000000000000000000000000000000000000; // D (0x0002004000000000) 
    12'h2c7 : errs =          63'b000000000000010000000001000000000000000000000000000000000000000; // D (0x0002008000000000) 
    12'ha5c : errs =          63'b000000000000010000000010000000000000000000000000000000000000000; // D (0x0002010000000000) 
    12'he53 : errs =          63'b000000000000010000000100000000000000000000000000000000000000000; // D (0x0002020000000000) 
    12'h64d : errs =          63'b000000000000010000001000000000000000000000000000000000000000000; // D (0x0002040000000000) 
    12'h348 : errs =          63'b000000000000010000010000000000000000000000000000000000000000000; // D (0x0002080000000000) 
    12'h942 : errs =          63'b000000000000010000100000000000000000000000000000000000000000000; // D (0x0002100000000000) 
    12'h86f : errs =          63'b000000000000010001000000000000000000000000000000000000000000000; // D (0x0002200000000000) 
    12'ha35 : errs =          63'b000000000000010010000000000000000000000000000000000000000000000; // D (0x0002400000000000) 
    12'he81 : errs =          63'b000000000000010100000000000000000000000000000000000000000000000; // D (0x0002800000000000) 
    12'h7e9 : errs =          63'b000000000000011000000000000000000000000000000000000000000000000; // D (0x0003000000000000) 
    12'h54e : errs =          63'b000000000000010000000000000000000000000000000000000000000000000; // S (0x0002000000000000) 
//    12'hfd2 : errs =          63'b000000000000110000000000000000000000000000000000000000000000000; // D (0x0006000000000000) 
//    12'h54f : errs =          63'b000000000001010000000000000000000000000000000000000000000000000; // D (0x000a000000000000) 
//    12'h54c : errs =          63'b000000000010010000000000000000000000000000000000000000000000000; // D (0x0012000000000000) 
//    12'h54a : errs =          63'b000000000100010000000000000000000000000000000000000000000000000; // D (0x0022000000000000) 
//    12'h546 : errs =          63'b000000001000010000000000000000000000000000000000000000000000000; // D (0x0042000000000000) 
//    12'h55e : errs =          63'b000000010000010000000000000000000000000000000000000000000000000; // D (0x0082000000000000) 
//    12'h56e : errs =          63'b000000100000010000000000000000000000000000000000000000000000000; // D (0x0102000000000000) 
//    12'h50e : errs =          63'b000001000000010000000000000000000000000000000000000000000000000; // D (0x0202000000000000) 
//    12'h5ce : errs =          63'b000010000000010000000000000000000000000000000000000000000000000; // D (0x0402000000000000) 
//    12'h44e : errs =          63'b000100000000010000000000000000000000000000000000000000000000000; // D (0x0802000000000000) 
//    12'h74e : errs =          63'b001000000000010000000000000000000000000000000000000000000000000; // D (0x1002000000000000) 
//    12'h14e : errs =          63'b010000000000010000000000000000000000000000000000000000000000000; // D (0x2002000000000000) 
//    12'hd4e : errs =          63'b100000000000010000000000000000000000000000000000000000000000000; // D (0x4002000000000000) 
    12'hfa5 : errs =          63'b000000000000100000000000000000000000000000000000000000000000001; // D (0x0004000000000001) 
    12'h0ee : errs =          63'b000000000000100000000000000000000000000000000000000000000000010; // D (0x0004000000000002) 
    12'hb41 : errs =          63'b000000000000100000000000000000000000000000000000000000000000100; // D (0x0004000000000004) 
    12'h926 : errs =          63'b000000000000100000000000000000000000000000000000000000000001000; // D (0x0004000000000008) 
    12'hde8 : errs =          63'b000000000000100000000000000000000000000000000000000000000010000; // D (0x0004000000000010) 
    12'h474 : errs =          63'b000000000000100000000000000000000000000000000000000000000100000; // D (0x0004000000000020) 
    12'h275 : errs =          63'b000000000000100000000000000000000000000000000000000000001000000; // D (0x0004000000000040) 
    12'he77 : errs =          63'b000000000000100000000000000000000000000000000000000000010000000; // D (0x0004000000000080) 
    12'h34a : errs =          63'b000000000000100000000000000000000000000000000000000000100000000; // D (0x0004000000000100) 
    12'hc09 : errs =          63'b000000000000100000000000000000000000000000000000000001000000000; // D (0x0004000000000200) 
    12'h7b6 : errs =          63'b000000000000100000000000000000000000000000000000000010000000000; // D (0x0004000000000400) 
    12'h5f1 : errs =          63'b000000000000100000000000000000000000000000000000000100000000000; // D (0x0004000000000800) 
    12'h17f : errs =          63'b000000000000100000000000000000000000000000000000001000000000000; // D (0x0004000000001000) 
    12'h863 : errs =          63'b000000000000100000000000000000000000000000000000010000000000000; // D (0x0004000000002000) 
    12'hf62 : errs =          63'b000000000000100000000000000000000000000000000000100000000000000; // D (0x0004000000004000) 
    12'h160 : errs =          63'b000000000000100000000000000000000000000000000001000000000000000; // D (0x0004000000008000) 
    12'h85d : errs =          63'b000000000000100000000000000000000000000000000010000000000000000; // D (0x0004000000010000) 
    12'hf1e : errs =          63'b000000000000100000000000000000000000000000000100000000000000000; // D (0x0004000000020000) 
    12'h198 : errs =          63'b000000000000100000000000000000000000000000001000000000000000000; // D (0x0004000000040000) 
    12'h9ad : errs =          63'b000000000000100000000000000000000000000000010000000000000000000; // D (0x0004000000080000) 
    12'hcfe : errs =          63'b000000000000100000000000000000000000000000100000000000000000000; // D (0x0004000000100000) 
    12'h658 : errs =          63'b000000000000100000000000000000000000000001000000000000000000000; // D (0x0004000000200000) 
    12'h62d : errs =          63'b000000000000100000000000000000000000000010000000000000000000000; // D (0x0004000000400000) 
    12'h6c7 : errs =          63'b000000000000100000000000000000000000000100000000000000000000000; // D (0x0004000000800000) 
    12'h713 : errs =          63'b000000000000100000000000000000000000001000000000000000000000000; // D (0x0004000001000000) 
    12'h4bb : errs =          63'b000000000000100000000000000000000000010000000000000000000000000; // D (0x0004000002000000) 
    12'h3eb : errs =          63'b000000000000100000000000000000000000100000000000000000000000000; // D (0x0004000004000000) 
    12'hd4b : errs =          63'b000000000000100000000000000000000001000000000000000000000000000; // D (0x0004000008000000) 
    12'h532 : errs =          63'b000000000000100000000000000000000010000000000000000000000000000; // D (0x0004000010000000) 
    12'h0f9 : errs =          63'b000000000000100000000000000000000100000000000000000000000000000; // D (0x0004000020000000) 
    12'hb6f : errs =          63'b000000000000100000000000000000001000000000000000000000000000000; // D (0x0004000040000000) 
    12'h97a : errs =          63'b000000000000100000000000000000010000000000000000000000000000000; // D (0x0004000080000000) 
    12'hd50 : errs =          63'b000000000000100000000000000000100000000000000000000000000000000; // D (0x0004000100000000) 
    12'h504 : errs =          63'b000000000000100000000000000001000000000000000000000000000000000; // D (0x0004000200000000) 
    12'h095 : errs =          63'b000000000000100000000000000010000000000000000000000000000000000; // D (0x0004000400000000) 
    12'hbb7 : errs =          63'b000000000000100000000000000100000000000000000000000000000000000; // D (0x0004000800000000) 
    12'h8ca : errs =          63'b000000000000100000000000001000000000000000000000000000000000000; // D (0x0004001000000000) 
    12'he30 : errs =          63'b000000000000100000000000010000000000000000000000000000000000000; // D (0x0004002000000000) 
    12'h3c4 : errs =          63'b000000000000100000000000100000000000000000000000000000000000000; // D (0x0004004000000000) 
    12'hd15 : errs =          63'b000000000000100000000001000000000000000000000000000000000000000; // D (0x0004008000000000) 
    12'h58e : errs =          63'b000000000000100000000010000000000000000000000000000000000000000; // D (0x0004010000000000) 
    12'h181 : errs =          63'b000000000000100000000100000000000000000000000000000000000000000; // D (0x0004020000000000) 
    12'h99f : errs =          63'b000000000000100000001000000000000000000000000000000000000000000; // D (0x0004040000000000) 
    12'hc9a : errs =          63'b000000000000100000010000000000000000000000000000000000000000000; // D (0x0004080000000000) 
    12'h690 : errs =          63'b000000000000100000100000000000000000000000000000000000000000000; // D (0x0004100000000000) 
    12'h7bd : errs =          63'b000000000000100001000000000000000000000000000000000000000000000; // D (0x0004200000000000) 
    12'h5e7 : errs =          63'b000000000000100010000000000000000000000000000000000000000000000; // D (0x0004400000000000) 
    12'h153 : errs =          63'b000000000000100100000000000000000000000000000000000000000000000; // D (0x0004800000000000) 
    12'h83b : errs =          63'b000000000000101000000000000000000000000000000000000000000000000; // D (0x0005000000000000) 
    12'hfd2 : errs =          63'b000000000000110000000000000000000000000000000000000000000000000; // D (0x0006000000000000) 
    12'ha9c : errs =          63'b000000000000100000000000000000000000000000000000000000000000000; // S (0x0004000000000000) 
//    12'ha9d : errs =          63'b000000000001100000000000000000000000000000000000000000000000000; // D (0x000c000000000000) 
//    12'ha9e : errs =          63'b000000000010100000000000000000000000000000000000000000000000000; // D (0x0014000000000000) 
//    12'ha98 : errs =          63'b000000000100100000000000000000000000000000000000000000000000000; // D (0x0024000000000000) 
//    12'ha94 : errs =          63'b000000001000100000000000000000000000000000000000000000000000000; // D (0x0044000000000000) 
//    12'ha8c : errs =          63'b000000010000100000000000000000000000000000000000000000000000000; // D (0x0084000000000000) 
//    12'habc : errs =          63'b000000100000100000000000000000000000000000000000000000000000000; // D (0x0104000000000000) 
//    12'hadc : errs =          63'b000001000000100000000000000000000000000000000000000000000000000; // D (0x0204000000000000) 
//    12'ha1c : errs =          63'b000010000000100000000000000000000000000000000000000000000000000; // D (0x0404000000000000) 
//    12'hb9c : errs =          63'b000100000000100000000000000000000000000000000000000000000000000; // D (0x0804000000000000) 
//    12'h89c : errs =          63'b001000000000100000000000000000000000000000000000000000000000000; // D (0x1004000000000000) 
//    12'he9c : errs =          63'b010000000000100000000000000000000000000000000000000000000000000; // D (0x2004000000000000) 
//    12'h29c : errs =          63'b100000000000100000000000000000000000000000000000000000000000000; // D (0x4004000000000000) 
    12'h538 : errs =          63'b000000000001000000000000000000000000000000000000000000000000001; // D (0x0008000000000001) 
    12'ha73 : errs =          63'b000000000001000000000000000000000000000000000000000000000000010; // D (0x0008000000000002) 
    12'h1dc : errs =          63'b000000000001000000000000000000000000000000000000000000000000100; // D (0x0008000000000004) 
    12'h3bb : errs =          63'b000000000001000000000000000000000000000000000000000000000001000; // D (0x0008000000000008) 
    12'h775 : errs =          63'b000000000001000000000000000000000000000000000000000000000010000; // D (0x0008000000000010) 
    12'hee9 : errs =          63'b000000000001000000000000000000000000000000000000000000000100000; // D (0x0008000000000020) 
    12'h8e8 : errs =          63'b000000000001000000000000000000000000000000000000000000001000000; // D (0x0008000000000040) 
    12'h4ea : errs =          63'b000000000001000000000000000000000000000000000000000000010000000; // D (0x0008000000000080) 
    12'h9d7 : errs =          63'b000000000001000000000000000000000000000000000000000000100000000; // D (0x0008000000000100) 
    12'h694 : errs =          63'b000000000001000000000000000000000000000000000000000001000000000; // D (0x0008000000000200) 
    12'hd2b : errs =          63'b000000000001000000000000000000000000000000000000000010000000000; // D (0x0008000000000400) 
    12'hf6c : errs =          63'b000000000001000000000000000000000000000000000000000100000000000; // D (0x0008000000000800) 
    12'hbe2 : errs =          63'b000000000001000000000000000000000000000000000000001000000000000; // D (0x0008000000001000) 
    12'h2fe : errs =          63'b000000000001000000000000000000000000000000000000010000000000000; // D (0x0008000000002000) 
    12'h5ff : errs =          63'b000000000001000000000000000000000000000000000000100000000000000; // D (0x0008000000004000) 
    12'hbfd : errs =          63'b000000000001000000000000000000000000000000000001000000000000000; // D (0x0008000000008000) 
    12'h2c0 : errs =          63'b000000000001000000000000000000000000000000000010000000000000000; // D (0x0008000000010000) 
    12'h583 : errs =          63'b000000000001000000000000000000000000000000000100000000000000000; // D (0x0008000000020000) 
    12'hb05 : errs =          63'b000000000001000000000000000000000000000000001000000000000000000; // D (0x0008000000040000) 
    12'h330 : errs =          63'b000000000001000000000000000000000000000000010000000000000000000; // D (0x0008000000080000) 
    12'h663 : errs =          63'b000000000001000000000000000000000000000000100000000000000000000; // D (0x0008000000100000) 
    12'hcc5 : errs =          63'b000000000001000000000000000000000000000001000000000000000000000; // D (0x0008000000200000) 
    12'hcb0 : errs =          63'b000000000001000000000000000000000000000010000000000000000000000; // D (0x0008000000400000) 
    12'hc5a : errs =          63'b000000000001000000000000000000000000000100000000000000000000000; // D (0x0008000000800000) 
    12'hd8e : errs =          63'b000000000001000000000000000000000000001000000000000000000000000; // D (0x0008000001000000) 
    12'he26 : errs =          63'b000000000001000000000000000000000000010000000000000000000000000; // D (0x0008000002000000) 
    12'h976 : errs =          63'b000000000001000000000000000000000000100000000000000000000000000; // D (0x0008000004000000) 
    12'h7d6 : errs =          63'b000000000001000000000000000000000001000000000000000000000000000; // D (0x0008000008000000) 
    12'hfaf : errs =          63'b000000000001000000000000000000000010000000000000000000000000000; // D (0x0008000010000000) 
    12'ha64 : errs =          63'b000000000001000000000000000000000100000000000000000000000000000; // D (0x0008000020000000) 
    12'h1f2 : errs =          63'b000000000001000000000000000000001000000000000000000000000000000; // D (0x0008000040000000) 
    12'h3e7 : errs =          63'b000000000001000000000000000000010000000000000000000000000000000; // D (0x0008000080000000) 
    12'h7cd : errs =          63'b000000000001000000000000000000100000000000000000000000000000000; // D (0x0008000100000000) 
    12'hf99 : errs =          63'b000000000001000000000000000001000000000000000000000000000000000; // D (0x0008000200000000) 
    12'ha08 : errs =          63'b000000000001000000000000000010000000000000000000000000000000000; // D (0x0008000400000000) 
    12'h12a : errs =          63'b000000000001000000000000000100000000000000000000000000000000000; // D (0x0008000800000000) 
    12'h257 : errs =          63'b000000000001000000000000001000000000000000000000000000000000000; // D (0x0008001000000000) 
    12'h4ad : errs =          63'b000000000001000000000000010000000000000000000000000000000000000; // D (0x0008002000000000) 
    12'h959 : errs =          63'b000000000001000000000000100000000000000000000000000000000000000; // D (0x0008004000000000) 
    12'h788 : errs =          63'b000000000001000000000001000000000000000000000000000000000000000; // D (0x0008008000000000) 
    12'hf13 : errs =          63'b000000000001000000000010000000000000000000000000000000000000000; // D (0x0008010000000000) 
    12'hb1c : errs =          63'b000000000001000000000100000000000000000000000000000000000000000; // D (0x0008020000000000) 
    12'h302 : errs =          63'b000000000001000000001000000000000000000000000000000000000000000; // D (0x0008040000000000) 
    12'h607 : errs =          63'b000000000001000000010000000000000000000000000000000000000000000; // D (0x0008080000000000) 
    12'hc0d : errs =          63'b000000000001000000100000000000000000000000000000000000000000000; // D (0x0008100000000000) 
    12'hd20 : errs =          63'b000000000001000001000000000000000000000000000000000000000000000; // D (0x0008200000000000) 
    12'hf7a : errs =          63'b000000000001000010000000000000000000000000000000000000000000000; // D (0x0008400000000000) 
    12'hbce : errs =          63'b000000000001000100000000000000000000000000000000000000000000000; // D (0x0008800000000000) 
    12'h2a6 : errs =          63'b000000000001001000000000000000000000000000000000000000000000000; // D (0x0009000000000000) 
    12'h54f : errs =          63'b000000000001010000000000000000000000000000000000000000000000000; // D (0x000a000000000000) 
    12'ha9d : errs =          63'b000000000001100000000000000000000000000000000000000000000000000; // D (0x000c000000000000) 
    12'h001 : errs =          63'b000000000001000000000000000000000000000000000000000000000000000; // S (0x0008000000000000) 
//    12'h003 : errs =          63'b000000000011000000000000000000000000000000000000000000000000000; // D (0x0018000000000000) 
//    12'h005 : errs =          63'b000000000101000000000000000000000000000000000000000000000000000; // D (0x0028000000000000) 
//    12'h009 : errs =          63'b000000001001000000000000000000000000000000000000000000000000000; // D (0x0048000000000000) 
//    12'h011 : errs =          63'b000000010001000000000000000000000000000000000000000000000000000; // D (0x0088000000000000) 
//    12'h021 : errs =          63'b000000100001000000000000000000000000000000000000000000000000000; // D (0x0108000000000000) 
//    12'h041 : errs =          63'b000001000001000000000000000000000000000000000000000000000000000; // D (0x0208000000000000) 
//    12'h081 : errs =          63'b000010000001000000000000000000000000000000000000000000000000000; // D (0x0408000000000000) 
//    12'h101 : errs =          63'b000100000001000000000000000000000000000000000000000000000000000; // D (0x0808000000000000) 
//    12'h201 : errs =          63'b001000000001000000000000000000000000000000000000000000000000000; // D (0x1008000000000000) 
//    12'h401 : errs =          63'b010000000001000000000000000000000000000000000000000000000000000; // D (0x2008000000000000) 
//    12'h801 : errs =          63'b100000000001000000000000000000000000000000000000000000000000000; // D (0x4008000000000000) 
    12'h53b : errs =          63'b000000000010000000000000000000000000000000000000000000000000001; // D (0x0010000000000001) 
    12'ha70 : errs =          63'b000000000010000000000000000000000000000000000000000000000000010; // D (0x0010000000000002) 
    12'h1df : errs =          63'b000000000010000000000000000000000000000000000000000000000000100; // D (0x0010000000000004) 
    12'h3b8 : errs =          63'b000000000010000000000000000000000000000000000000000000000001000; // D (0x0010000000000008) 
    12'h776 : errs =          63'b000000000010000000000000000000000000000000000000000000000010000; // D (0x0010000000000010) 
    12'heea : errs =          63'b000000000010000000000000000000000000000000000000000000000100000; // D (0x0010000000000020) 
    12'h8eb : errs =          63'b000000000010000000000000000000000000000000000000000000001000000; // D (0x0010000000000040) 
    12'h4e9 : errs =          63'b000000000010000000000000000000000000000000000000000000010000000; // D (0x0010000000000080) 
    12'h9d4 : errs =          63'b000000000010000000000000000000000000000000000000000000100000000; // D (0x0010000000000100) 
    12'h697 : errs =          63'b000000000010000000000000000000000000000000000000000001000000000; // D (0x0010000000000200) 
    12'hd28 : errs =          63'b000000000010000000000000000000000000000000000000000010000000000; // D (0x0010000000000400) 
    12'hf6f : errs =          63'b000000000010000000000000000000000000000000000000000100000000000; // D (0x0010000000000800) 
    12'hbe1 : errs =          63'b000000000010000000000000000000000000000000000000001000000000000; // D (0x0010000000001000) 
    12'h2fd : errs =          63'b000000000010000000000000000000000000000000000000010000000000000; // D (0x0010000000002000) 
    12'h5fc : errs =          63'b000000000010000000000000000000000000000000000000100000000000000; // D (0x0010000000004000) 
    12'hbfe : errs =          63'b000000000010000000000000000000000000000000000001000000000000000; // D (0x0010000000008000) 
    12'h2c3 : errs =          63'b000000000010000000000000000000000000000000000010000000000000000; // D (0x0010000000010000) 
    12'h580 : errs =          63'b000000000010000000000000000000000000000000000100000000000000000; // D (0x0010000000020000) 
    12'hb06 : errs =          63'b000000000010000000000000000000000000000000001000000000000000000; // D (0x0010000000040000) 
    12'h333 : errs =          63'b000000000010000000000000000000000000000000010000000000000000000; // D (0x0010000000080000) 
    12'h660 : errs =          63'b000000000010000000000000000000000000000000100000000000000000000; // D (0x0010000000100000) 
    12'hcc6 : errs =          63'b000000000010000000000000000000000000000001000000000000000000000; // D (0x0010000000200000) 
    12'hcb3 : errs =          63'b000000000010000000000000000000000000000010000000000000000000000; // D (0x0010000000400000) 
    12'hc59 : errs =          63'b000000000010000000000000000000000000000100000000000000000000000; // D (0x0010000000800000) 
    12'hd8d : errs =          63'b000000000010000000000000000000000000001000000000000000000000000; // D (0x0010000001000000) 
    12'he25 : errs =          63'b000000000010000000000000000000000000010000000000000000000000000; // D (0x0010000002000000) 
    12'h975 : errs =          63'b000000000010000000000000000000000000100000000000000000000000000; // D (0x0010000004000000) 
    12'h7d5 : errs =          63'b000000000010000000000000000000000001000000000000000000000000000; // D (0x0010000008000000) 
    12'hfac : errs =          63'b000000000010000000000000000000000010000000000000000000000000000; // D (0x0010000010000000) 
    12'ha67 : errs =          63'b000000000010000000000000000000000100000000000000000000000000000; // D (0x0010000020000000) 
    12'h1f1 : errs =          63'b000000000010000000000000000000001000000000000000000000000000000; // D (0x0010000040000000) 
    12'h3e4 : errs =          63'b000000000010000000000000000000010000000000000000000000000000000; // D (0x0010000080000000) 
    12'h7ce : errs =          63'b000000000010000000000000000000100000000000000000000000000000000; // D (0x0010000100000000) 
    12'hf9a : errs =          63'b000000000010000000000000000001000000000000000000000000000000000; // D (0x0010000200000000) 
    12'ha0b : errs =          63'b000000000010000000000000000010000000000000000000000000000000000; // D (0x0010000400000000) 
    12'h129 : errs =          63'b000000000010000000000000000100000000000000000000000000000000000; // D (0x0010000800000000) 
    12'h254 : errs =          63'b000000000010000000000000001000000000000000000000000000000000000; // D (0x0010001000000000) 
    12'h4ae : errs =          63'b000000000010000000000000010000000000000000000000000000000000000; // D (0x0010002000000000) 
    12'h95a : errs =          63'b000000000010000000000000100000000000000000000000000000000000000; // D (0x0010004000000000) 
    12'h78b : errs =          63'b000000000010000000000001000000000000000000000000000000000000000; // D (0x0010008000000000) 
    12'hf10 : errs =          63'b000000000010000000000010000000000000000000000000000000000000000; // D (0x0010010000000000) 
    12'hb1f : errs =          63'b000000000010000000000100000000000000000000000000000000000000000; // D (0x0010020000000000) 
    12'h301 : errs =          63'b000000000010000000001000000000000000000000000000000000000000000; // D (0x0010040000000000) 
    12'h604 : errs =          63'b000000000010000000010000000000000000000000000000000000000000000; // D (0x0010080000000000) 
    12'hc0e : errs =          63'b000000000010000000100000000000000000000000000000000000000000000; // D (0x0010100000000000) 
    12'hd23 : errs =          63'b000000000010000001000000000000000000000000000000000000000000000; // D (0x0010200000000000) 
    12'hf79 : errs =          63'b000000000010000010000000000000000000000000000000000000000000000; // D (0x0010400000000000) 
    12'hbcd : errs =          63'b000000000010000100000000000000000000000000000000000000000000000; // D (0x0010800000000000) 
    12'h2a5 : errs =          63'b000000000010001000000000000000000000000000000000000000000000000; // D (0x0011000000000000) 
    12'h54c : errs =          63'b000000000010010000000000000000000000000000000000000000000000000; // D (0x0012000000000000) 
    12'ha9e : errs =          63'b000000000010100000000000000000000000000000000000000000000000000; // D (0x0014000000000000) 
    12'h003 : errs =          63'b000000000011000000000000000000000000000000000000000000000000000; // D (0x0018000000000000) 
    12'h002 : errs =          63'b000000000010000000000000000000000000000000000000000000000000000; // S (0x0010000000000000) 
//    12'h006 : errs =          63'b000000000110000000000000000000000000000000000000000000000000000; // D (0x0030000000000000) 
//    12'h00a : errs =          63'b000000001010000000000000000000000000000000000000000000000000000; // D (0x0050000000000000) 
//    12'h012 : errs =          63'b000000010010000000000000000000000000000000000000000000000000000; // D (0x0090000000000000) 
//    12'h022 : errs =          63'b000000100010000000000000000000000000000000000000000000000000000; // D (0x0110000000000000) 
//    12'h042 : errs =          63'b000001000010000000000000000000000000000000000000000000000000000; // D (0x0210000000000000) 
//    12'h082 : errs =          63'b000010000010000000000000000000000000000000000000000000000000000; // D (0x0410000000000000) 
//    12'h102 : errs =          63'b000100000010000000000000000000000000000000000000000000000000000; // D (0x0810000000000000) 
//    12'h202 : errs =          63'b001000000010000000000000000000000000000000000000000000000000000; // D (0x1010000000000000) 
//    12'h402 : errs =          63'b010000000010000000000000000000000000000000000000000000000000000; // D (0x2010000000000000) 
//    12'h802 : errs =          63'b100000000010000000000000000000000000000000000000000000000000000; // D (0x4010000000000000) 
    12'h53d : errs =          63'b000000000100000000000000000000000000000000000000000000000000001; // D (0x0020000000000001) 
    12'ha76 : errs =          63'b000000000100000000000000000000000000000000000000000000000000010; // D (0x0020000000000002) 
    12'h1d9 : errs =          63'b000000000100000000000000000000000000000000000000000000000000100; // D (0x0020000000000004) 
    12'h3be : errs =          63'b000000000100000000000000000000000000000000000000000000000001000; // D (0x0020000000000008) 
    12'h770 : errs =          63'b000000000100000000000000000000000000000000000000000000000010000; // D (0x0020000000000010) 
    12'heec : errs =          63'b000000000100000000000000000000000000000000000000000000000100000; // D (0x0020000000000020) 
    12'h8ed : errs =          63'b000000000100000000000000000000000000000000000000000000001000000; // D (0x0020000000000040) 
    12'h4ef : errs =          63'b000000000100000000000000000000000000000000000000000000010000000; // D (0x0020000000000080) 
    12'h9d2 : errs =          63'b000000000100000000000000000000000000000000000000000000100000000; // D (0x0020000000000100) 
    12'h691 : errs =          63'b000000000100000000000000000000000000000000000000000001000000000; // D (0x0020000000000200) 
    12'hd2e : errs =          63'b000000000100000000000000000000000000000000000000000010000000000; // D (0x0020000000000400) 
    12'hf69 : errs =          63'b000000000100000000000000000000000000000000000000000100000000000; // D (0x0020000000000800) 
    12'hbe7 : errs =          63'b000000000100000000000000000000000000000000000000001000000000000; // D (0x0020000000001000) 
    12'h2fb : errs =          63'b000000000100000000000000000000000000000000000000010000000000000; // D (0x0020000000002000) 
    12'h5fa : errs =          63'b000000000100000000000000000000000000000000000000100000000000000; // D (0x0020000000004000) 
    12'hbf8 : errs =          63'b000000000100000000000000000000000000000000000001000000000000000; // D (0x0020000000008000) 
    12'h2c5 : errs =          63'b000000000100000000000000000000000000000000000010000000000000000; // D (0x0020000000010000) 
    12'h586 : errs =          63'b000000000100000000000000000000000000000000000100000000000000000; // D (0x0020000000020000) 
    12'hb00 : errs =          63'b000000000100000000000000000000000000000000001000000000000000000; // D (0x0020000000040000) 
    12'h335 : errs =          63'b000000000100000000000000000000000000000000010000000000000000000; // D (0x0020000000080000) 
    12'h666 : errs =          63'b000000000100000000000000000000000000000000100000000000000000000; // D (0x0020000000100000) 
    12'hcc0 : errs =          63'b000000000100000000000000000000000000000001000000000000000000000; // D (0x0020000000200000) 
    12'hcb5 : errs =          63'b000000000100000000000000000000000000000010000000000000000000000; // D (0x0020000000400000) 
    12'hc5f : errs =          63'b000000000100000000000000000000000000000100000000000000000000000; // D (0x0020000000800000) 
    12'hd8b : errs =          63'b000000000100000000000000000000000000001000000000000000000000000; // D (0x0020000001000000) 
    12'he23 : errs =          63'b000000000100000000000000000000000000010000000000000000000000000; // D (0x0020000002000000) 
    12'h973 : errs =          63'b000000000100000000000000000000000000100000000000000000000000000; // D (0x0020000004000000) 
    12'h7d3 : errs =          63'b000000000100000000000000000000000001000000000000000000000000000; // D (0x0020000008000000) 
    12'hfaa : errs =          63'b000000000100000000000000000000000010000000000000000000000000000; // D (0x0020000010000000) 
    12'ha61 : errs =          63'b000000000100000000000000000000000100000000000000000000000000000; // D (0x0020000020000000) 
    12'h1f7 : errs =          63'b000000000100000000000000000000001000000000000000000000000000000; // D (0x0020000040000000) 
    12'h3e2 : errs =          63'b000000000100000000000000000000010000000000000000000000000000000; // D (0x0020000080000000) 
    12'h7c8 : errs =          63'b000000000100000000000000000000100000000000000000000000000000000; // D (0x0020000100000000) 
    12'hf9c : errs =          63'b000000000100000000000000000001000000000000000000000000000000000; // D (0x0020000200000000) 
    12'ha0d : errs =          63'b000000000100000000000000000010000000000000000000000000000000000; // D (0x0020000400000000) 
    12'h12f : errs =          63'b000000000100000000000000000100000000000000000000000000000000000; // D (0x0020000800000000) 
    12'h252 : errs =          63'b000000000100000000000000001000000000000000000000000000000000000; // D (0x0020001000000000) 
    12'h4a8 : errs =          63'b000000000100000000000000010000000000000000000000000000000000000; // D (0x0020002000000000) 
    12'h95c : errs =          63'b000000000100000000000000100000000000000000000000000000000000000; // D (0x0020004000000000) 
    12'h78d : errs =          63'b000000000100000000000001000000000000000000000000000000000000000; // D (0x0020008000000000) 
    12'hf16 : errs =          63'b000000000100000000000010000000000000000000000000000000000000000; // D (0x0020010000000000) 
    12'hb19 : errs =          63'b000000000100000000000100000000000000000000000000000000000000000; // D (0x0020020000000000) 
    12'h307 : errs =          63'b000000000100000000001000000000000000000000000000000000000000000; // D (0x0020040000000000) 
    12'h602 : errs =          63'b000000000100000000010000000000000000000000000000000000000000000; // D (0x0020080000000000) 
    12'hc08 : errs =          63'b000000000100000000100000000000000000000000000000000000000000000; // D (0x0020100000000000) 
    12'hd25 : errs =          63'b000000000100000001000000000000000000000000000000000000000000000; // D (0x0020200000000000) 
    12'hf7f : errs =          63'b000000000100000010000000000000000000000000000000000000000000000; // D (0x0020400000000000) 
    12'hbcb : errs =          63'b000000000100000100000000000000000000000000000000000000000000000; // D (0x0020800000000000) 
    12'h2a3 : errs =          63'b000000000100001000000000000000000000000000000000000000000000000; // D (0x0021000000000000) 
    12'h54a : errs =          63'b000000000100010000000000000000000000000000000000000000000000000; // D (0x0022000000000000) 
    12'ha98 : errs =          63'b000000000100100000000000000000000000000000000000000000000000000; // D (0x0024000000000000) 
    12'h005 : errs =          63'b000000000101000000000000000000000000000000000000000000000000000; // D (0x0028000000000000) 
    12'h006 : errs =          63'b000000000110000000000000000000000000000000000000000000000000000; // D (0x0030000000000000) 
    12'h004 : errs =          63'b000000000100000000000000000000000000000000000000000000000000000; // S (0x0020000000000000) 
//    12'h00c : errs =          63'b000000001100000000000000000000000000000000000000000000000000000; // D (0x0060000000000000) 
//    12'h014 : errs =          63'b000000010100000000000000000000000000000000000000000000000000000; // D (0x00a0000000000000) 
//    12'h024 : errs =          63'b000000100100000000000000000000000000000000000000000000000000000; // D (0x0120000000000000) 
//    12'h044 : errs =          63'b000001000100000000000000000000000000000000000000000000000000000; // D (0x0220000000000000) 
//    12'h084 : errs =          63'b000010000100000000000000000000000000000000000000000000000000000; // D (0x0420000000000000) 
//    12'h104 : errs =          63'b000100000100000000000000000000000000000000000000000000000000000; // D (0x0820000000000000) 
//    12'h204 : errs =          63'b001000000100000000000000000000000000000000000000000000000000000; // D (0x1020000000000000) 
//    12'h404 : errs =          63'b010000000100000000000000000000000000000000000000000000000000000; // D (0x2020000000000000) 
//    12'h804 : errs =          63'b100000000100000000000000000000000000000000000000000000000000000; // D (0x4020000000000000) 
    12'h531 : errs =          63'b000000001000000000000000000000000000000000000000000000000000001; // D (0x0040000000000001) 
    12'ha7a : errs =          63'b000000001000000000000000000000000000000000000000000000000000010; // D (0x0040000000000002) 
    12'h1d5 : errs =          63'b000000001000000000000000000000000000000000000000000000000000100; // D (0x0040000000000004) 
    12'h3b2 : errs =          63'b000000001000000000000000000000000000000000000000000000000001000; // D (0x0040000000000008) 
    12'h77c : errs =          63'b000000001000000000000000000000000000000000000000000000000010000; // D (0x0040000000000010) 
    12'hee0 : errs =          63'b000000001000000000000000000000000000000000000000000000000100000; // D (0x0040000000000020) 
    12'h8e1 : errs =          63'b000000001000000000000000000000000000000000000000000000001000000; // D (0x0040000000000040) 
    12'h4e3 : errs =          63'b000000001000000000000000000000000000000000000000000000010000000; // D (0x0040000000000080) 
    12'h9de : errs =          63'b000000001000000000000000000000000000000000000000000000100000000; // D (0x0040000000000100) 
    12'h69d : errs =          63'b000000001000000000000000000000000000000000000000000001000000000; // D (0x0040000000000200) 
    12'hd22 : errs =          63'b000000001000000000000000000000000000000000000000000010000000000; // D (0x0040000000000400) 
    12'hf65 : errs =          63'b000000001000000000000000000000000000000000000000000100000000000; // D (0x0040000000000800) 
    12'hbeb : errs =          63'b000000001000000000000000000000000000000000000000001000000000000; // D (0x0040000000001000) 
    12'h2f7 : errs =          63'b000000001000000000000000000000000000000000000000010000000000000; // D (0x0040000000002000) 
    12'h5f6 : errs =          63'b000000001000000000000000000000000000000000000000100000000000000; // D (0x0040000000004000) 
    12'hbf4 : errs =          63'b000000001000000000000000000000000000000000000001000000000000000; // D (0x0040000000008000) 
    12'h2c9 : errs =          63'b000000001000000000000000000000000000000000000010000000000000000; // D (0x0040000000010000) 
    12'h58a : errs =          63'b000000001000000000000000000000000000000000000100000000000000000; // D (0x0040000000020000) 
    12'hb0c : errs =          63'b000000001000000000000000000000000000000000001000000000000000000; // D (0x0040000000040000) 
    12'h339 : errs =          63'b000000001000000000000000000000000000000000010000000000000000000; // D (0x0040000000080000) 
    12'h66a : errs =          63'b000000001000000000000000000000000000000000100000000000000000000; // D (0x0040000000100000) 
    12'hccc : errs =          63'b000000001000000000000000000000000000000001000000000000000000000; // D (0x0040000000200000) 
    12'hcb9 : errs =          63'b000000001000000000000000000000000000000010000000000000000000000; // D (0x0040000000400000) 
    12'hc53 : errs =          63'b000000001000000000000000000000000000000100000000000000000000000; // D (0x0040000000800000) 
    12'hd87 : errs =          63'b000000001000000000000000000000000000001000000000000000000000000; // D (0x0040000001000000) 
    12'he2f : errs =          63'b000000001000000000000000000000000000010000000000000000000000000; // D (0x0040000002000000) 
    12'h97f : errs =          63'b000000001000000000000000000000000000100000000000000000000000000; // D (0x0040000004000000) 
    12'h7df : errs =          63'b000000001000000000000000000000000001000000000000000000000000000; // D (0x0040000008000000) 
    12'hfa6 : errs =          63'b000000001000000000000000000000000010000000000000000000000000000; // D (0x0040000010000000) 
    12'ha6d : errs =          63'b000000001000000000000000000000000100000000000000000000000000000; // D (0x0040000020000000) 
    12'h1fb : errs =          63'b000000001000000000000000000000001000000000000000000000000000000; // D (0x0040000040000000) 
    12'h3ee : errs =          63'b000000001000000000000000000000010000000000000000000000000000000; // D (0x0040000080000000) 
    12'h7c4 : errs =          63'b000000001000000000000000000000100000000000000000000000000000000; // D (0x0040000100000000) 
    12'hf90 : errs =          63'b000000001000000000000000000001000000000000000000000000000000000; // D (0x0040000200000000) 
    12'ha01 : errs =          63'b000000001000000000000000000010000000000000000000000000000000000; // D (0x0040000400000000) 
    12'h123 : errs =          63'b000000001000000000000000000100000000000000000000000000000000000; // D (0x0040000800000000) 
    12'h25e : errs =          63'b000000001000000000000000001000000000000000000000000000000000000; // D (0x0040001000000000) 
    12'h4a4 : errs =          63'b000000001000000000000000010000000000000000000000000000000000000; // D (0x0040002000000000) 
    12'h950 : errs =          63'b000000001000000000000000100000000000000000000000000000000000000; // D (0x0040004000000000) 
    12'h781 : errs =          63'b000000001000000000000001000000000000000000000000000000000000000; // D (0x0040008000000000) 
    12'hf1a : errs =          63'b000000001000000000000010000000000000000000000000000000000000000; // D (0x0040010000000000) 
    12'hb15 : errs =          63'b000000001000000000000100000000000000000000000000000000000000000; // D (0x0040020000000000) 
    12'h30b : errs =          63'b000000001000000000001000000000000000000000000000000000000000000; // D (0x0040040000000000) 
    12'h60e : errs =          63'b000000001000000000010000000000000000000000000000000000000000000; // D (0x0040080000000000) 
    12'hc04 : errs =          63'b000000001000000000100000000000000000000000000000000000000000000; // D (0x0040100000000000) 
    12'hd29 : errs =          63'b000000001000000001000000000000000000000000000000000000000000000; // D (0x0040200000000000) 
    12'hf73 : errs =          63'b000000001000000010000000000000000000000000000000000000000000000; // D (0x0040400000000000) 
    12'hbc7 : errs =          63'b000000001000000100000000000000000000000000000000000000000000000; // D (0x0040800000000000) 
    12'h2af : errs =          63'b000000001000001000000000000000000000000000000000000000000000000; // D (0x0041000000000000) 
    12'h546 : errs =          63'b000000001000010000000000000000000000000000000000000000000000000; // D (0x0042000000000000) 
    12'ha94 : errs =          63'b000000001000100000000000000000000000000000000000000000000000000; // D (0x0044000000000000) 
    12'h009 : errs =          63'b000000001001000000000000000000000000000000000000000000000000000; // D (0x0048000000000000) 
    12'h00a : errs =          63'b000000001010000000000000000000000000000000000000000000000000000; // D (0x0050000000000000) 
    12'h00c : errs =          63'b000000001100000000000000000000000000000000000000000000000000000; // D (0x0060000000000000) 
    12'h008 : errs =          63'b000000001000000000000000000000000000000000000000000000000000000; // S (0x0040000000000000) 
//    12'h018 : errs =          63'b000000011000000000000000000000000000000000000000000000000000000; // D (0x00c0000000000000) 
//    12'h028 : errs =          63'b000000101000000000000000000000000000000000000000000000000000000; // D (0x0140000000000000) 
//    12'h048 : errs =          63'b000001001000000000000000000000000000000000000000000000000000000; // D (0x0240000000000000) 
//    12'h088 : errs =          63'b000010001000000000000000000000000000000000000000000000000000000; // D (0x0440000000000000) 
//    12'h108 : errs =          63'b000100001000000000000000000000000000000000000000000000000000000; // D (0x0840000000000000) 
//    12'h208 : errs =          63'b001000001000000000000000000000000000000000000000000000000000000; // D (0x1040000000000000) 
//    12'h408 : errs =          63'b010000001000000000000000000000000000000000000000000000000000000; // D (0x2040000000000000) 
//    12'h808 : errs =          63'b100000001000000000000000000000000000000000000000000000000000000; // D (0x4040000000000000) 
    12'h529 : errs =          63'b000000010000000000000000000000000000000000000000000000000000001; // D (0x0080000000000001) 
    12'ha62 : errs =          63'b000000010000000000000000000000000000000000000000000000000000010; // D (0x0080000000000002) 
    12'h1cd : errs =          63'b000000010000000000000000000000000000000000000000000000000000100; // D (0x0080000000000004) 
    12'h3aa : errs =          63'b000000010000000000000000000000000000000000000000000000000001000; // D (0x0080000000000008) 
    12'h764 : errs =          63'b000000010000000000000000000000000000000000000000000000000010000; // D (0x0080000000000010) 
    12'hef8 : errs =          63'b000000010000000000000000000000000000000000000000000000000100000; // D (0x0080000000000020) 
    12'h8f9 : errs =          63'b000000010000000000000000000000000000000000000000000000001000000; // D (0x0080000000000040) 
    12'h4fb : errs =          63'b000000010000000000000000000000000000000000000000000000010000000; // D (0x0080000000000080) 
    12'h9c6 : errs =          63'b000000010000000000000000000000000000000000000000000000100000000; // D (0x0080000000000100) 
    12'h685 : errs =          63'b000000010000000000000000000000000000000000000000000001000000000; // D (0x0080000000000200) 
    12'hd3a : errs =          63'b000000010000000000000000000000000000000000000000000010000000000; // D (0x0080000000000400) 
    12'hf7d : errs =          63'b000000010000000000000000000000000000000000000000000100000000000; // D (0x0080000000000800) 
    12'hbf3 : errs =          63'b000000010000000000000000000000000000000000000000001000000000000; // D (0x0080000000001000) 
    12'h2ef : errs =          63'b000000010000000000000000000000000000000000000000010000000000000; // D (0x0080000000002000) 
    12'h5ee : errs =          63'b000000010000000000000000000000000000000000000000100000000000000; // D (0x0080000000004000) 
    12'hbec : errs =          63'b000000010000000000000000000000000000000000000001000000000000000; // D (0x0080000000008000) 
    12'h2d1 : errs =          63'b000000010000000000000000000000000000000000000010000000000000000; // D (0x0080000000010000) 
    12'h592 : errs =          63'b000000010000000000000000000000000000000000000100000000000000000; // D (0x0080000000020000) 
    12'hb14 : errs =          63'b000000010000000000000000000000000000000000001000000000000000000; // D (0x0080000000040000) 
    12'h321 : errs =          63'b000000010000000000000000000000000000000000010000000000000000000; // D (0x0080000000080000) 
    12'h672 : errs =          63'b000000010000000000000000000000000000000000100000000000000000000; // D (0x0080000000100000) 
    12'hcd4 : errs =          63'b000000010000000000000000000000000000000001000000000000000000000; // D (0x0080000000200000) 
    12'hca1 : errs =          63'b000000010000000000000000000000000000000010000000000000000000000; // D (0x0080000000400000) 
    12'hc4b : errs =          63'b000000010000000000000000000000000000000100000000000000000000000; // D (0x0080000000800000) 
    12'hd9f : errs =          63'b000000010000000000000000000000000000001000000000000000000000000; // D (0x0080000001000000) 
    12'he37 : errs =          63'b000000010000000000000000000000000000010000000000000000000000000; // D (0x0080000002000000) 
    12'h967 : errs =          63'b000000010000000000000000000000000000100000000000000000000000000; // D (0x0080000004000000) 
    12'h7c7 : errs =          63'b000000010000000000000000000000000001000000000000000000000000000; // D (0x0080000008000000) 
    12'hfbe : errs =          63'b000000010000000000000000000000000010000000000000000000000000000; // D (0x0080000010000000) 
    12'ha75 : errs =          63'b000000010000000000000000000000000100000000000000000000000000000; // D (0x0080000020000000) 
    12'h1e3 : errs =          63'b000000010000000000000000000000001000000000000000000000000000000; // D (0x0080000040000000) 
    12'h3f6 : errs =          63'b000000010000000000000000000000010000000000000000000000000000000; // D (0x0080000080000000) 
    12'h7dc : errs =          63'b000000010000000000000000000000100000000000000000000000000000000; // D (0x0080000100000000) 
    12'hf88 : errs =          63'b000000010000000000000000000001000000000000000000000000000000000; // D (0x0080000200000000) 
    12'ha19 : errs =          63'b000000010000000000000000000010000000000000000000000000000000000; // D (0x0080000400000000) 
    12'h13b : errs =          63'b000000010000000000000000000100000000000000000000000000000000000; // D (0x0080000800000000) 
    12'h246 : errs =          63'b000000010000000000000000001000000000000000000000000000000000000; // D (0x0080001000000000) 
    12'h4bc : errs =          63'b000000010000000000000000010000000000000000000000000000000000000; // D (0x0080002000000000) 
    12'h948 : errs =          63'b000000010000000000000000100000000000000000000000000000000000000; // D (0x0080004000000000) 
    12'h799 : errs =          63'b000000010000000000000001000000000000000000000000000000000000000; // D (0x0080008000000000) 
    12'hf02 : errs =          63'b000000010000000000000010000000000000000000000000000000000000000; // D (0x0080010000000000) 
    12'hb0d : errs =          63'b000000010000000000000100000000000000000000000000000000000000000; // D (0x0080020000000000) 
    12'h313 : errs =          63'b000000010000000000001000000000000000000000000000000000000000000; // D (0x0080040000000000) 
    12'h616 : errs =          63'b000000010000000000010000000000000000000000000000000000000000000; // D (0x0080080000000000) 
    12'hc1c : errs =          63'b000000010000000000100000000000000000000000000000000000000000000; // D (0x0080100000000000) 
    12'hd31 : errs =          63'b000000010000000001000000000000000000000000000000000000000000000; // D (0x0080200000000000) 
    12'hf6b : errs =          63'b000000010000000010000000000000000000000000000000000000000000000; // D (0x0080400000000000) 
    12'hbdf : errs =          63'b000000010000000100000000000000000000000000000000000000000000000; // D (0x0080800000000000) 
    12'h2b7 : errs =          63'b000000010000001000000000000000000000000000000000000000000000000; // D (0x0081000000000000) 
    12'h55e : errs =          63'b000000010000010000000000000000000000000000000000000000000000000; // D (0x0082000000000000) 
    12'ha8c : errs =          63'b000000010000100000000000000000000000000000000000000000000000000; // D (0x0084000000000000) 
    12'h011 : errs =          63'b000000010001000000000000000000000000000000000000000000000000000; // D (0x0088000000000000) 
    12'h012 : errs =          63'b000000010010000000000000000000000000000000000000000000000000000; // D (0x0090000000000000) 
    12'h014 : errs =          63'b000000010100000000000000000000000000000000000000000000000000000; // D (0x00a0000000000000) 
    12'h018 : errs =          63'b000000011000000000000000000000000000000000000000000000000000000; // D (0x00c0000000000000) 
    12'h010 : errs =          63'b000000010000000000000000000000000000000000000000000000000000000; // S (0x0080000000000000) 
//    12'h030 : errs =          63'b000000110000000000000000000000000000000000000000000000000000000; // D (0x0180000000000000) 
//    12'h050 : errs =          63'b000001010000000000000000000000000000000000000000000000000000000; // D (0x0280000000000000) 
//    12'h090 : errs =          63'b000010010000000000000000000000000000000000000000000000000000000; // D (0x0480000000000000) 
//    12'h110 : errs =          63'b000100010000000000000000000000000000000000000000000000000000000; // D (0x0880000000000000) 
//    12'h210 : errs =          63'b001000010000000000000000000000000000000000000000000000000000000; // D (0x1080000000000000) 
//    12'h410 : errs =          63'b010000010000000000000000000000000000000000000000000000000000000; // D (0x2080000000000000) 
//    12'h810 : errs =          63'b100000010000000000000000000000000000000000000000000000000000000; // D (0x4080000000000000) 
    12'h519 : errs =          63'b000000100000000000000000000000000000000000000000000000000000001; // D (0x0100000000000001) 
    12'ha52 : errs =          63'b000000100000000000000000000000000000000000000000000000000000010; // D (0x0100000000000002) 
    12'h1fd : errs =          63'b000000100000000000000000000000000000000000000000000000000000100; // D (0x0100000000000004) 
    12'h39a : errs =          63'b000000100000000000000000000000000000000000000000000000000001000; // D (0x0100000000000008) 
    12'h754 : errs =          63'b000000100000000000000000000000000000000000000000000000000010000; // D (0x0100000000000010) 
    12'hec8 : errs =          63'b000000100000000000000000000000000000000000000000000000000100000; // D (0x0100000000000020) 
    12'h8c9 : errs =          63'b000000100000000000000000000000000000000000000000000000001000000; // D (0x0100000000000040) 
    12'h4cb : errs =          63'b000000100000000000000000000000000000000000000000000000010000000; // D (0x0100000000000080) 
    12'h9f6 : errs =          63'b000000100000000000000000000000000000000000000000000000100000000; // D (0x0100000000000100) 
    12'h6b5 : errs =          63'b000000100000000000000000000000000000000000000000000001000000000; // D (0x0100000000000200) 
    12'hd0a : errs =          63'b000000100000000000000000000000000000000000000000000010000000000; // D (0x0100000000000400) 
    12'hf4d : errs =          63'b000000100000000000000000000000000000000000000000000100000000000; // D (0x0100000000000800) 
    12'hbc3 : errs =          63'b000000100000000000000000000000000000000000000000001000000000000; // D (0x0100000000001000) 
    12'h2df : errs =          63'b000000100000000000000000000000000000000000000000010000000000000; // D (0x0100000000002000) 
    12'h5de : errs =          63'b000000100000000000000000000000000000000000000000100000000000000; // D (0x0100000000004000) 
    12'hbdc : errs =          63'b000000100000000000000000000000000000000000000001000000000000000; // D (0x0100000000008000) 
    12'h2e1 : errs =          63'b000000100000000000000000000000000000000000000010000000000000000; // D (0x0100000000010000) 
    12'h5a2 : errs =          63'b000000100000000000000000000000000000000000000100000000000000000; // D (0x0100000000020000) 
    12'hb24 : errs =          63'b000000100000000000000000000000000000000000001000000000000000000; // D (0x0100000000040000) 
    12'h311 : errs =          63'b000000100000000000000000000000000000000000010000000000000000000; // D (0x0100000000080000) 
    12'h642 : errs =          63'b000000100000000000000000000000000000000000100000000000000000000; // D (0x0100000000100000) 
    12'hce4 : errs =          63'b000000100000000000000000000000000000000001000000000000000000000; // D (0x0100000000200000) 
    12'hc91 : errs =          63'b000000100000000000000000000000000000000010000000000000000000000; // D (0x0100000000400000) 
    12'hc7b : errs =          63'b000000100000000000000000000000000000000100000000000000000000000; // D (0x0100000000800000) 
    12'hdaf : errs =          63'b000000100000000000000000000000000000001000000000000000000000000; // D (0x0100000001000000) 
    12'he07 : errs =          63'b000000100000000000000000000000000000010000000000000000000000000; // D (0x0100000002000000) 
    12'h957 : errs =          63'b000000100000000000000000000000000000100000000000000000000000000; // D (0x0100000004000000) 
    12'h7f7 : errs =          63'b000000100000000000000000000000000001000000000000000000000000000; // D (0x0100000008000000) 
    12'hf8e : errs =          63'b000000100000000000000000000000000010000000000000000000000000000; // D (0x0100000010000000) 
    12'ha45 : errs =          63'b000000100000000000000000000000000100000000000000000000000000000; // D (0x0100000020000000) 
    12'h1d3 : errs =          63'b000000100000000000000000000000001000000000000000000000000000000; // D (0x0100000040000000) 
    12'h3c6 : errs =          63'b000000100000000000000000000000010000000000000000000000000000000; // D (0x0100000080000000) 
    12'h7ec : errs =          63'b000000100000000000000000000000100000000000000000000000000000000; // D (0x0100000100000000) 
    12'hfb8 : errs =          63'b000000100000000000000000000001000000000000000000000000000000000; // D (0x0100000200000000) 
    12'ha29 : errs =          63'b000000100000000000000000000010000000000000000000000000000000000; // D (0x0100000400000000) 
    12'h10b : errs =          63'b000000100000000000000000000100000000000000000000000000000000000; // D (0x0100000800000000) 
    12'h276 : errs =          63'b000000100000000000000000001000000000000000000000000000000000000; // D (0x0100001000000000) 
    12'h48c : errs =          63'b000000100000000000000000010000000000000000000000000000000000000; // D (0x0100002000000000) 
    12'h978 : errs =          63'b000000100000000000000000100000000000000000000000000000000000000; // D (0x0100004000000000) 
    12'h7a9 : errs =          63'b000000100000000000000001000000000000000000000000000000000000000; // D (0x0100008000000000) 
    12'hf32 : errs =          63'b000000100000000000000010000000000000000000000000000000000000000; // D (0x0100010000000000) 
    12'hb3d : errs =          63'b000000100000000000000100000000000000000000000000000000000000000; // D (0x0100020000000000) 
    12'h323 : errs =          63'b000000100000000000001000000000000000000000000000000000000000000; // D (0x0100040000000000) 
    12'h626 : errs =          63'b000000100000000000010000000000000000000000000000000000000000000; // D (0x0100080000000000) 
    12'hc2c : errs =          63'b000000100000000000100000000000000000000000000000000000000000000; // D (0x0100100000000000) 
    12'hd01 : errs =          63'b000000100000000001000000000000000000000000000000000000000000000; // D (0x0100200000000000) 
    12'hf5b : errs =          63'b000000100000000010000000000000000000000000000000000000000000000; // D (0x0100400000000000) 
    12'hbef : errs =          63'b000000100000000100000000000000000000000000000000000000000000000; // D (0x0100800000000000) 
    12'h287 : errs =          63'b000000100000001000000000000000000000000000000000000000000000000; // D (0x0101000000000000) 
    12'h56e : errs =          63'b000000100000010000000000000000000000000000000000000000000000000; // D (0x0102000000000000) 
    12'habc : errs =          63'b000000100000100000000000000000000000000000000000000000000000000; // D (0x0104000000000000) 
    12'h021 : errs =          63'b000000100001000000000000000000000000000000000000000000000000000; // D (0x0108000000000000) 
    12'h022 : errs =          63'b000000100010000000000000000000000000000000000000000000000000000; // D (0x0110000000000000) 
    12'h024 : errs =          63'b000000100100000000000000000000000000000000000000000000000000000; // D (0x0120000000000000) 
    12'h028 : errs =          63'b000000101000000000000000000000000000000000000000000000000000000; // D (0x0140000000000000) 
    12'h030 : errs =          63'b000000110000000000000000000000000000000000000000000000000000000; // D (0x0180000000000000) 
    12'h020 : errs =          63'b000000100000000000000000000000000000000000000000000000000000000; // S (0x0100000000000000) 
//    12'h060 : errs =          63'b000001100000000000000000000000000000000000000000000000000000000; // D (0x0300000000000000) 
//    12'h0a0 : errs =          63'b000010100000000000000000000000000000000000000000000000000000000; // D (0x0500000000000000) 
//    12'h120 : errs =          63'b000100100000000000000000000000000000000000000000000000000000000; // D (0x0900000000000000) 
//    12'h220 : errs =          63'b001000100000000000000000000000000000000000000000000000000000000; // D (0x1100000000000000) 
//    12'h420 : errs =          63'b010000100000000000000000000000000000000000000000000000000000000; // D (0x2100000000000000) 
//    12'h820 : errs =          63'b100000100000000000000000000000000000000000000000000000000000000; // D (0x4100000000000000) 
    12'h579 : errs =          63'b000001000000000000000000000000000000000000000000000000000000001; // D (0x0200000000000001) 
    12'ha32 : errs =          63'b000001000000000000000000000000000000000000000000000000000000010; // D (0x0200000000000002) 
    12'h19d : errs =          63'b000001000000000000000000000000000000000000000000000000000000100; // D (0x0200000000000004) 
    12'h3fa : errs =          63'b000001000000000000000000000000000000000000000000000000000001000; // D (0x0200000000000008) 
    12'h734 : errs =          63'b000001000000000000000000000000000000000000000000000000000010000; // D (0x0200000000000010) 
    12'hea8 : errs =          63'b000001000000000000000000000000000000000000000000000000000100000; // D (0x0200000000000020) 
    12'h8a9 : errs =          63'b000001000000000000000000000000000000000000000000000000001000000; // D (0x0200000000000040) 
    12'h4ab : errs =          63'b000001000000000000000000000000000000000000000000000000010000000; // D (0x0200000000000080) 
    12'h996 : errs =          63'b000001000000000000000000000000000000000000000000000000100000000; // D (0x0200000000000100) 
    12'h6d5 : errs =          63'b000001000000000000000000000000000000000000000000000001000000000; // D (0x0200000000000200) 
    12'hd6a : errs =          63'b000001000000000000000000000000000000000000000000000010000000000; // D (0x0200000000000400) 
    12'hf2d : errs =          63'b000001000000000000000000000000000000000000000000000100000000000; // D (0x0200000000000800) 
    12'hba3 : errs =          63'b000001000000000000000000000000000000000000000000001000000000000; // D (0x0200000000001000) 
    12'h2bf : errs =          63'b000001000000000000000000000000000000000000000000010000000000000; // D (0x0200000000002000) 
    12'h5be : errs =          63'b000001000000000000000000000000000000000000000000100000000000000; // D (0x0200000000004000) 
    12'hbbc : errs =          63'b000001000000000000000000000000000000000000000001000000000000000; // D (0x0200000000008000) 
    12'h281 : errs =          63'b000001000000000000000000000000000000000000000010000000000000000; // D (0x0200000000010000) 
    12'h5c2 : errs =          63'b000001000000000000000000000000000000000000000100000000000000000; // D (0x0200000000020000) 
    12'hb44 : errs =          63'b000001000000000000000000000000000000000000001000000000000000000; // D (0x0200000000040000) 
    12'h371 : errs =          63'b000001000000000000000000000000000000000000010000000000000000000; // D (0x0200000000080000) 
    12'h622 : errs =          63'b000001000000000000000000000000000000000000100000000000000000000; // D (0x0200000000100000) 
    12'hc84 : errs =          63'b000001000000000000000000000000000000000001000000000000000000000; // D (0x0200000000200000) 
    12'hcf1 : errs =          63'b000001000000000000000000000000000000000010000000000000000000000; // D (0x0200000000400000) 
    12'hc1b : errs =          63'b000001000000000000000000000000000000000100000000000000000000000; // D (0x0200000000800000) 
    12'hdcf : errs =          63'b000001000000000000000000000000000000001000000000000000000000000; // D (0x0200000001000000) 
    12'he67 : errs =          63'b000001000000000000000000000000000000010000000000000000000000000; // D (0x0200000002000000) 
    12'h937 : errs =          63'b000001000000000000000000000000000000100000000000000000000000000; // D (0x0200000004000000) 
    12'h797 : errs =          63'b000001000000000000000000000000000001000000000000000000000000000; // D (0x0200000008000000) 
    12'hfee : errs =          63'b000001000000000000000000000000000010000000000000000000000000000; // D (0x0200000010000000) 
    12'ha25 : errs =          63'b000001000000000000000000000000000100000000000000000000000000000; // D (0x0200000020000000) 
    12'h1b3 : errs =          63'b000001000000000000000000000000001000000000000000000000000000000; // D (0x0200000040000000) 
    12'h3a6 : errs =          63'b000001000000000000000000000000010000000000000000000000000000000; // D (0x0200000080000000) 
    12'h78c : errs =          63'b000001000000000000000000000000100000000000000000000000000000000; // D (0x0200000100000000) 
    12'hfd8 : errs =          63'b000001000000000000000000000001000000000000000000000000000000000; // D (0x0200000200000000) 
    12'ha49 : errs =          63'b000001000000000000000000000010000000000000000000000000000000000; // D (0x0200000400000000) 
    12'h16b : errs =          63'b000001000000000000000000000100000000000000000000000000000000000; // D (0x0200000800000000) 
    12'h216 : errs =          63'b000001000000000000000000001000000000000000000000000000000000000; // D (0x0200001000000000) 
    12'h4ec : errs =          63'b000001000000000000000000010000000000000000000000000000000000000; // D (0x0200002000000000) 
    12'h918 : errs =          63'b000001000000000000000000100000000000000000000000000000000000000; // D (0x0200004000000000) 
    12'h7c9 : errs =          63'b000001000000000000000001000000000000000000000000000000000000000; // D (0x0200008000000000) 
    12'hf52 : errs =          63'b000001000000000000000010000000000000000000000000000000000000000; // D (0x0200010000000000) 
    12'hb5d : errs =          63'b000001000000000000000100000000000000000000000000000000000000000; // D (0x0200020000000000) 
    12'h343 : errs =          63'b000001000000000000001000000000000000000000000000000000000000000; // D (0x0200040000000000) 
    12'h646 : errs =          63'b000001000000000000010000000000000000000000000000000000000000000; // D (0x0200080000000000) 
    12'hc4c : errs =          63'b000001000000000000100000000000000000000000000000000000000000000; // D (0x0200100000000000) 
    12'hd61 : errs =          63'b000001000000000001000000000000000000000000000000000000000000000; // D (0x0200200000000000) 
    12'hf3b : errs =          63'b000001000000000010000000000000000000000000000000000000000000000; // D (0x0200400000000000) 
    12'hb8f : errs =          63'b000001000000000100000000000000000000000000000000000000000000000; // D (0x0200800000000000) 
    12'h2e7 : errs =          63'b000001000000001000000000000000000000000000000000000000000000000; // D (0x0201000000000000) 
    12'h50e : errs =          63'b000001000000010000000000000000000000000000000000000000000000000; // D (0x0202000000000000) 
    12'hadc : errs =          63'b000001000000100000000000000000000000000000000000000000000000000; // D (0x0204000000000000) 
    12'h041 : errs =          63'b000001000001000000000000000000000000000000000000000000000000000; // D (0x0208000000000000) 
    12'h042 : errs =          63'b000001000010000000000000000000000000000000000000000000000000000; // D (0x0210000000000000) 
    12'h044 : errs =          63'b000001000100000000000000000000000000000000000000000000000000000; // D (0x0220000000000000) 
    12'h048 : errs =          63'b000001001000000000000000000000000000000000000000000000000000000; // D (0x0240000000000000) 
    12'h050 : errs =          63'b000001010000000000000000000000000000000000000000000000000000000; // D (0x0280000000000000) 
    12'h060 : errs =          63'b000001100000000000000000000000000000000000000000000000000000000; // D (0x0300000000000000) 
    12'h040 : errs =          63'b000001000000000000000000000000000000000000000000000000000000000; // S (0x0200000000000000) 
//    12'h0c0 : errs =          63'b000011000000000000000000000000000000000000000000000000000000000; // D (0x0600000000000000) 
//    12'h140 : errs =          63'b000101000000000000000000000000000000000000000000000000000000000; // D (0x0a00000000000000) 
//    12'h240 : errs =          63'b001001000000000000000000000000000000000000000000000000000000000; // D (0x1200000000000000) 
//    12'h440 : errs =          63'b010001000000000000000000000000000000000000000000000000000000000; // D (0x2200000000000000) 
//    12'h840 : errs =          63'b100001000000000000000000000000000000000000000000000000000000000; // D (0x4200000000000000) 
    12'h5b9 : errs =          63'b000010000000000000000000000000000000000000000000000000000000001; // D (0x0400000000000001) 
    12'haf2 : errs =          63'b000010000000000000000000000000000000000000000000000000000000010; // D (0x0400000000000002) 
    12'h15d : errs =          63'b000010000000000000000000000000000000000000000000000000000000100; // D (0x0400000000000004) 
    12'h33a : errs =          63'b000010000000000000000000000000000000000000000000000000000001000; // D (0x0400000000000008) 
    12'h7f4 : errs =          63'b000010000000000000000000000000000000000000000000000000000010000; // D (0x0400000000000010) 
    12'he68 : errs =          63'b000010000000000000000000000000000000000000000000000000000100000; // D (0x0400000000000020) 
    12'h869 : errs =          63'b000010000000000000000000000000000000000000000000000000001000000; // D (0x0400000000000040) 
    12'h46b : errs =          63'b000010000000000000000000000000000000000000000000000000010000000; // D (0x0400000000000080) 
    12'h956 : errs =          63'b000010000000000000000000000000000000000000000000000000100000000; // D (0x0400000000000100) 
    12'h615 : errs =          63'b000010000000000000000000000000000000000000000000000001000000000; // D (0x0400000000000200) 
    12'hdaa : errs =          63'b000010000000000000000000000000000000000000000000000010000000000; // D (0x0400000000000400) 
    12'hfed : errs =          63'b000010000000000000000000000000000000000000000000000100000000000; // D (0x0400000000000800) 
    12'hb63 : errs =          63'b000010000000000000000000000000000000000000000000001000000000000; // D (0x0400000000001000) 
    12'h27f : errs =          63'b000010000000000000000000000000000000000000000000010000000000000; // D (0x0400000000002000) 
    12'h57e : errs =          63'b000010000000000000000000000000000000000000000000100000000000000; // D (0x0400000000004000) 
    12'hb7c : errs =          63'b000010000000000000000000000000000000000000000001000000000000000; // D (0x0400000000008000) 
    12'h241 : errs =          63'b000010000000000000000000000000000000000000000010000000000000000; // D (0x0400000000010000) 
    12'h502 : errs =          63'b000010000000000000000000000000000000000000000100000000000000000; // D (0x0400000000020000) 
    12'hb84 : errs =          63'b000010000000000000000000000000000000000000001000000000000000000; // D (0x0400000000040000) 
    12'h3b1 : errs =          63'b000010000000000000000000000000000000000000010000000000000000000; // D (0x0400000000080000) 
    12'h6e2 : errs =          63'b000010000000000000000000000000000000000000100000000000000000000; // D (0x0400000000100000) 
    12'hc44 : errs =          63'b000010000000000000000000000000000000000001000000000000000000000; // D (0x0400000000200000) 
    12'hc31 : errs =          63'b000010000000000000000000000000000000000010000000000000000000000; // D (0x0400000000400000) 
    12'hcdb : errs =          63'b000010000000000000000000000000000000000100000000000000000000000; // D (0x0400000000800000) 
    12'hd0f : errs =          63'b000010000000000000000000000000000000001000000000000000000000000; // D (0x0400000001000000) 
    12'hea7 : errs =          63'b000010000000000000000000000000000000010000000000000000000000000; // D (0x0400000002000000) 
    12'h9f7 : errs =          63'b000010000000000000000000000000000000100000000000000000000000000; // D (0x0400000004000000) 
    12'h757 : errs =          63'b000010000000000000000000000000000001000000000000000000000000000; // D (0x0400000008000000) 
    12'hf2e : errs =          63'b000010000000000000000000000000000010000000000000000000000000000; // D (0x0400000010000000) 
    12'hae5 : errs =          63'b000010000000000000000000000000000100000000000000000000000000000; // D (0x0400000020000000) 
    12'h173 : errs =          63'b000010000000000000000000000000001000000000000000000000000000000; // D (0x0400000040000000) 
    12'h366 : errs =          63'b000010000000000000000000000000010000000000000000000000000000000; // D (0x0400000080000000) 
    12'h74c : errs =          63'b000010000000000000000000000000100000000000000000000000000000000; // D (0x0400000100000000) 
    12'hf18 : errs =          63'b000010000000000000000000000001000000000000000000000000000000000; // D (0x0400000200000000) 
    12'ha89 : errs =          63'b000010000000000000000000000010000000000000000000000000000000000; // D (0x0400000400000000) 
    12'h1ab : errs =          63'b000010000000000000000000000100000000000000000000000000000000000; // D (0x0400000800000000) 
    12'h2d6 : errs =          63'b000010000000000000000000001000000000000000000000000000000000000; // D (0x0400001000000000) 
    12'h42c : errs =          63'b000010000000000000000000010000000000000000000000000000000000000; // D (0x0400002000000000) 
    12'h9d8 : errs =          63'b000010000000000000000000100000000000000000000000000000000000000; // D (0x0400004000000000) 
    12'h709 : errs =          63'b000010000000000000000001000000000000000000000000000000000000000; // D (0x0400008000000000) 
    12'hf92 : errs =          63'b000010000000000000000010000000000000000000000000000000000000000; // D (0x0400010000000000) 
    12'hb9d : errs =          63'b000010000000000000000100000000000000000000000000000000000000000; // D (0x0400020000000000) 
    12'h383 : errs =          63'b000010000000000000001000000000000000000000000000000000000000000; // D (0x0400040000000000) 
    12'h686 : errs =          63'b000010000000000000010000000000000000000000000000000000000000000; // D (0x0400080000000000) 
    12'hc8c : errs =          63'b000010000000000000100000000000000000000000000000000000000000000; // D (0x0400100000000000) 
    12'hda1 : errs =          63'b000010000000000001000000000000000000000000000000000000000000000; // D (0x0400200000000000) 
    12'hffb : errs =          63'b000010000000000010000000000000000000000000000000000000000000000; // D (0x0400400000000000) 
    12'hb4f : errs =          63'b000010000000000100000000000000000000000000000000000000000000000; // D (0x0400800000000000) 
    12'h227 : errs =          63'b000010000000001000000000000000000000000000000000000000000000000; // D (0x0401000000000000) 
    12'h5ce : errs =          63'b000010000000010000000000000000000000000000000000000000000000000; // D (0x0402000000000000) 
    12'ha1c : errs =          63'b000010000000100000000000000000000000000000000000000000000000000; // D (0x0404000000000000) 
    12'h081 : errs =          63'b000010000001000000000000000000000000000000000000000000000000000; // D (0x0408000000000000) 
    12'h082 : errs =          63'b000010000010000000000000000000000000000000000000000000000000000; // D (0x0410000000000000) 
    12'h084 : errs =          63'b000010000100000000000000000000000000000000000000000000000000000; // D (0x0420000000000000) 
    12'h088 : errs =          63'b000010001000000000000000000000000000000000000000000000000000000; // D (0x0440000000000000) 
    12'h090 : errs =          63'b000010010000000000000000000000000000000000000000000000000000000; // D (0x0480000000000000) 
    12'h0a0 : errs =          63'b000010100000000000000000000000000000000000000000000000000000000; // D (0x0500000000000000) 
    12'h0c0 : errs =          63'b000011000000000000000000000000000000000000000000000000000000000; // D (0x0600000000000000) 
    12'h080 : errs =          63'b000010000000000000000000000000000000000000000000000000000000000; // S (0x0400000000000000) 
//    12'h180 : errs =          63'b000110000000000000000000000000000000000000000000000000000000000; // D (0x0c00000000000000) 
//    12'h280 : errs =          63'b001010000000000000000000000000000000000000000000000000000000000; // D (0x1400000000000000) 
//    12'h480 : errs =          63'b010010000000000000000000000000000000000000000000000000000000000; // D (0x2400000000000000) 
//    12'h880 : errs =          63'b100010000000000000000000000000000000000000000000000000000000000; // D (0x4400000000000000) 
    12'h439 : errs =          63'b000100000000000000000000000000000000000000000000000000000000001; // D (0x0800000000000001) 
    12'hb72 : errs =          63'b000100000000000000000000000000000000000000000000000000000000010; // D (0x0800000000000002) 
    12'h0dd : errs =          63'b000100000000000000000000000000000000000000000000000000000000100; // D (0x0800000000000004) 
    12'h2ba : errs =          63'b000100000000000000000000000000000000000000000000000000000001000; // D (0x0800000000000008) 
    12'h674 : errs =          63'b000100000000000000000000000000000000000000000000000000000010000; // D (0x0800000000000010) 
    12'hfe8 : errs =          63'b000100000000000000000000000000000000000000000000000000000100000; // D (0x0800000000000020) 
    12'h9e9 : errs =          63'b000100000000000000000000000000000000000000000000000000001000000; // D (0x0800000000000040) 
    12'h5eb : errs =          63'b000100000000000000000000000000000000000000000000000000010000000; // D (0x0800000000000080) 
    12'h8d6 : errs =          63'b000100000000000000000000000000000000000000000000000000100000000; // D (0x0800000000000100) 
    12'h795 : errs =          63'b000100000000000000000000000000000000000000000000000001000000000; // D (0x0800000000000200) 
    12'hc2a : errs =          63'b000100000000000000000000000000000000000000000000000010000000000; // D (0x0800000000000400) 
    12'he6d : errs =          63'b000100000000000000000000000000000000000000000000000100000000000; // D (0x0800000000000800) 
    12'hae3 : errs =          63'b000100000000000000000000000000000000000000000000001000000000000; // D (0x0800000000001000) 
    12'h3ff : errs =          63'b000100000000000000000000000000000000000000000000010000000000000; // D (0x0800000000002000) 
    12'h4fe : errs =          63'b000100000000000000000000000000000000000000000000100000000000000; // D (0x0800000000004000) 
    12'hafc : errs =          63'b000100000000000000000000000000000000000000000001000000000000000; // D (0x0800000000008000) 
    12'h3c1 : errs =          63'b000100000000000000000000000000000000000000000010000000000000000; // D (0x0800000000010000) 
    12'h482 : errs =          63'b000100000000000000000000000000000000000000000100000000000000000; // D (0x0800000000020000) 
    12'ha04 : errs =          63'b000100000000000000000000000000000000000000001000000000000000000; // D (0x0800000000040000) 
    12'h231 : errs =          63'b000100000000000000000000000000000000000000010000000000000000000; // D (0x0800000000080000) 
    12'h762 : errs =          63'b000100000000000000000000000000000000000000100000000000000000000; // D (0x0800000000100000) 
    12'hdc4 : errs =          63'b000100000000000000000000000000000000000001000000000000000000000; // D (0x0800000000200000) 
    12'hdb1 : errs =          63'b000100000000000000000000000000000000000010000000000000000000000; // D (0x0800000000400000) 
    12'hd5b : errs =          63'b000100000000000000000000000000000000000100000000000000000000000; // D (0x0800000000800000) 
    12'hc8f : errs =          63'b000100000000000000000000000000000000001000000000000000000000000; // D (0x0800000001000000) 
    12'hf27 : errs =          63'b000100000000000000000000000000000000010000000000000000000000000; // D (0x0800000002000000) 
    12'h877 : errs =          63'b000100000000000000000000000000000000100000000000000000000000000; // D (0x0800000004000000) 
    12'h6d7 : errs =          63'b000100000000000000000000000000000001000000000000000000000000000; // D (0x0800000008000000) 
    12'heae : errs =          63'b000100000000000000000000000000000010000000000000000000000000000; // D (0x0800000010000000) 
    12'hb65 : errs =          63'b000100000000000000000000000000000100000000000000000000000000000; // D (0x0800000020000000) 
    12'h0f3 : errs =          63'b000100000000000000000000000000001000000000000000000000000000000; // D (0x0800000040000000) 
    12'h2e6 : errs =          63'b000100000000000000000000000000010000000000000000000000000000000; // D (0x0800000080000000) 
    12'h6cc : errs =          63'b000100000000000000000000000000100000000000000000000000000000000; // D (0x0800000100000000) 
    12'he98 : errs =          63'b000100000000000000000000000001000000000000000000000000000000000; // D (0x0800000200000000) 
    12'hb09 : errs =          63'b000100000000000000000000000010000000000000000000000000000000000; // D (0x0800000400000000) 
    12'h02b : errs =          63'b000100000000000000000000000100000000000000000000000000000000000; // D (0x0800000800000000) 
    12'h356 : errs =          63'b000100000000000000000000001000000000000000000000000000000000000; // D (0x0800001000000000) 
    12'h5ac : errs =          63'b000100000000000000000000010000000000000000000000000000000000000; // D (0x0800002000000000) 
    12'h858 : errs =          63'b000100000000000000000000100000000000000000000000000000000000000; // D (0x0800004000000000) 
    12'h689 : errs =          63'b000100000000000000000001000000000000000000000000000000000000000; // D (0x0800008000000000) 
    12'he12 : errs =          63'b000100000000000000000010000000000000000000000000000000000000000; // D (0x0800010000000000) 
    12'ha1d : errs =          63'b000100000000000000000100000000000000000000000000000000000000000; // D (0x0800020000000000) 
    12'h203 : errs =          63'b000100000000000000001000000000000000000000000000000000000000000; // D (0x0800040000000000) 
    12'h706 : errs =          63'b000100000000000000010000000000000000000000000000000000000000000; // D (0x0800080000000000) 
    12'hd0c : errs =          63'b000100000000000000100000000000000000000000000000000000000000000; // D (0x0800100000000000) 
    12'hc21 : errs =          63'b000100000000000001000000000000000000000000000000000000000000000; // D (0x0800200000000000) 
    12'he7b : errs =          63'b000100000000000010000000000000000000000000000000000000000000000; // D (0x0800400000000000) 
    12'hacf : errs =          63'b000100000000000100000000000000000000000000000000000000000000000; // D (0x0800800000000000) 
    12'h3a7 : errs =          63'b000100000000001000000000000000000000000000000000000000000000000; // D (0x0801000000000000) 
    12'h44e : errs =          63'b000100000000010000000000000000000000000000000000000000000000000; // D (0x0802000000000000) 
    12'hb9c : errs =          63'b000100000000100000000000000000000000000000000000000000000000000; // D (0x0804000000000000) 
    12'h101 : errs =          63'b000100000001000000000000000000000000000000000000000000000000000; // D (0x0808000000000000) 
    12'h102 : errs =          63'b000100000010000000000000000000000000000000000000000000000000000; // D (0x0810000000000000) 
    12'h104 : errs =          63'b000100000100000000000000000000000000000000000000000000000000000; // D (0x0820000000000000) 
    12'h108 : errs =          63'b000100001000000000000000000000000000000000000000000000000000000; // D (0x0840000000000000) 
    12'h110 : errs =          63'b000100010000000000000000000000000000000000000000000000000000000; // D (0x0880000000000000) 
    12'h120 : errs =          63'b000100100000000000000000000000000000000000000000000000000000000; // D (0x0900000000000000) 
    12'h140 : errs =          63'b000101000000000000000000000000000000000000000000000000000000000; // D (0x0a00000000000000) 
    12'h180 : errs =          63'b000110000000000000000000000000000000000000000000000000000000000; // D (0x0c00000000000000) 
    12'h100 : errs =          63'b000100000000000000000000000000000000000000000000000000000000000; // S (0x0800000000000000) 
//    12'h300 : errs =          63'b001100000000000000000000000000000000000000000000000000000000000; // D (0x1800000000000000) 
//    12'h500 : errs =          63'b010100000000000000000000000000000000000000000000000000000000000; // D (0x2800000000000000) 
//    12'h900 : errs =          63'b100100000000000000000000000000000000000000000000000000000000000; // D (0x4800000000000000) 
    12'h739 : errs =          63'b001000000000000000000000000000000000000000000000000000000000001; // D (0x1000000000000001) 
    12'h872 : errs =          63'b001000000000000000000000000000000000000000000000000000000000010; // D (0x1000000000000002) 
    12'h3dd : errs =          63'b001000000000000000000000000000000000000000000000000000000000100; // D (0x1000000000000004) 
    12'h1ba : errs =          63'b001000000000000000000000000000000000000000000000000000000001000; // D (0x1000000000000008) 
    12'h574 : errs =          63'b001000000000000000000000000000000000000000000000000000000010000; // D (0x1000000000000010) 
    12'hce8 : errs =          63'b001000000000000000000000000000000000000000000000000000000100000; // D (0x1000000000000020) 
    12'hae9 : errs =          63'b001000000000000000000000000000000000000000000000000000001000000; // D (0x1000000000000040) 
    12'h6eb : errs =          63'b001000000000000000000000000000000000000000000000000000010000000; // D (0x1000000000000080) 
    12'hbd6 : errs =          63'b001000000000000000000000000000000000000000000000000000100000000; // D (0x1000000000000100) 
    12'h495 : errs =          63'b001000000000000000000000000000000000000000000000000001000000000; // D (0x1000000000000200) 
    12'hf2a : errs =          63'b001000000000000000000000000000000000000000000000000010000000000; // D (0x1000000000000400) 
    12'hd6d : errs =          63'b001000000000000000000000000000000000000000000000000100000000000; // D (0x1000000000000800) 
    12'h9e3 : errs =          63'b001000000000000000000000000000000000000000000000001000000000000; // D (0x1000000000001000) 
    12'h0ff : errs =          63'b001000000000000000000000000000000000000000000000010000000000000; // D (0x1000000000002000) 
    12'h7fe : errs =          63'b001000000000000000000000000000000000000000000000100000000000000; // D (0x1000000000004000) 
    12'h9fc : errs =          63'b001000000000000000000000000000000000000000000001000000000000000; // D (0x1000000000008000) 
    12'h0c1 : errs =          63'b001000000000000000000000000000000000000000000010000000000000000; // D (0x1000000000010000) 
    12'h782 : errs =          63'b001000000000000000000000000000000000000000000100000000000000000; // D (0x1000000000020000) 
    12'h904 : errs =          63'b001000000000000000000000000000000000000000001000000000000000000; // D (0x1000000000040000) 
    12'h131 : errs =          63'b001000000000000000000000000000000000000000010000000000000000000; // D (0x1000000000080000) 
    12'h462 : errs =          63'b001000000000000000000000000000000000000000100000000000000000000; // D (0x1000000000100000) 
    12'hec4 : errs =          63'b001000000000000000000000000000000000000001000000000000000000000; // D (0x1000000000200000) 
    12'heb1 : errs =          63'b001000000000000000000000000000000000000010000000000000000000000; // D (0x1000000000400000) 
    12'he5b : errs =          63'b001000000000000000000000000000000000000100000000000000000000000; // D (0x1000000000800000) 
    12'hf8f : errs =          63'b001000000000000000000000000000000000001000000000000000000000000; // D (0x1000000001000000) 
    12'hc27 : errs =          63'b001000000000000000000000000000000000010000000000000000000000000; // D (0x1000000002000000) 
    12'hb77 : errs =          63'b001000000000000000000000000000000000100000000000000000000000000; // D (0x1000000004000000) 
    12'h5d7 : errs =          63'b001000000000000000000000000000000001000000000000000000000000000; // D (0x1000000008000000) 
    12'hdae : errs =          63'b001000000000000000000000000000000010000000000000000000000000000; // D (0x1000000010000000) 
    12'h865 : errs =          63'b001000000000000000000000000000000100000000000000000000000000000; // D (0x1000000020000000) 
    12'h3f3 : errs =          63'b001000000000000000000000000000001000000000000000000000000000000; // D (0x1000000040000000) 
    12'h1e6 : errs =          63'b001000000000000000000000000000010000000000000000000000000000000; // D (0x1000000080000000) 
    12'h5cc : errs =          63'b001000000000000000000000000000100000000000000000000000000000000; // D (0x1000000100000000) 
    12'hd98 : errs =          63'b001000000000000000000000000001000000000000000000000000000000000; // D (0x1000000200000000) 
    12'h809 : errs =          63'b001000000000000000000000000010000000000000000000000000000000000; // D (0x1000000400000000) 
    12'h32b : errs =          63'b001000000000000000000000000100000000000000000000000000000000000; // D (0x1000000800000000) 
    12'h056 : errs =          63'b001000000000000000000000001000000000000000000000000000000000000; // D (0x1000001000000000) 
    12'h6ac : errs =          63'b001000000000000000000000010000000000000000000000000000000000000; // D (0x1000002000000000) 
    12'hb58 : errs =          63'b001000000000000000000000100000000000000000000000000000000000000; // D (0x1000004000000000) 
    12'h589 : errs =          63'b001000000000000000000001000000000000000000000000000000000000000; // D (0x1000008000000000) 
    12'hd12 : errs =          63'b001000000000000000000010000000000000000000000000000000000000000; // D (0x1000010000000000) 
    12'h91d : errs =          63'b001000000000000000000100000000000000000000000000000000000000000; // D (0x1000020000000000) 
    12'h103 : errs =          63'b001000000000000000001000000000000000000000000000000000000000000; // D (0x1000040000000000) 
    12'h406 : errs =          63'b001000000000000000010000000000000000000000000000000000000000000; // D (0x1000080000000000) 
    12'he0c : errs =          63'b001000000000000000100000000000000000000000000000000000000000000; // D (0x1000100000000000) 
    12'hf21 : errs =          63'b001000000000000001000000000000000000000000000000000000000000000; // D (0x1000200000000000) 
    12'hd7b : errs =          63'b001000000000000010000000000000000000000000000000000000000000000; // D (0x1000400000000000) 
    12'h9cf : errs =          63'b001000000000000100000000000000000000000000000000000000000000000; // D (0x1000800000000000) 
    12'h0a7 : errs =          63'b001000000000001000000000000000000000000000000000000000000000000; // D (0x1001000000000000) 
    12'h74e : errs =          63'b001000000000010000000000000000000000000000000000000000000000000; // D (0x1002000000000000) 
    12'h89c : errs =          63'b001000000000100000000000000000000000000000000000000000000000000; // D (0x1004000000000000) 
    12'h201 : errs =          63'b001000000001000000000000000000000000000000000000000000000000000; // D (0x1008000000000000) 
    12'h202 : errs =          63'b001000000010000000000000000000000000000000000000000000000000000; // D (0x1010000000000000) 
    12'h204 : errs =          63'b001000000100000000000000000000000000000000000000000000000000000; // D (0x1020000000000000) 
    12'h208 : errs =          63'b001000001000000000000000000000000000000000000000000000000000000; // D (0x1040000000000000) 
    12'h210 : errs =          63'b001000010000000000000000000000000000000000000000000000000000000; // D (0x1080000000000000) 
    12'h220 : errs =          63'b001000100000000000000000000000000000000000000000000000000000000; // D (0x1100000000000000) 
    12'h240 : errs =          63'b001001000000000000000000000000000000000000000000000000000000000; // D (0x1200000000000000) 
    12'h280 : errs =          63'b001010000000000000000000000000000000000000000000000000000000000; // D (0x1400000000000000) 
    12'h300 : errs =          63'b001100000000000000000000000000000000000000000000000000000000000; // D (0x1800000000000000) 
    12'h200 : errs =          63'b001000000000000000000000000000000000000000000000000000000000000; // S (0x1000000000000000) 
//    12'h600 : errs =          63'b011000000000000000000000000000000000000000000000000000000000000; // D (0x3000000000000000) 
//    12'ha00 : errs =          63'b101000000000000000000000000000000000000000000000000000000000000; // D (0x5000000000000000) 
    12'h139 : errs =          63'b010000000000000000000000000000000000000000000000000000000000001; // D (0x2000000000000001) 
    12'he72 : errs =          63'b010000000000000000000000000000000000000000000000000000000000010; // D (0x2000000000000002) 
    12'h5dd : errs =          63'b010000000000000000000000000000000000000000000000000000000000100; // D (0x2000000000000004) 
    12'h7ba : errs =          63'b010000000000000000000000000000000000000000000000000000000001000; // D (0x2000000000000008) 
    12'h374 : errs =          63'b010000000000000000000000000000000000000000000000000000000010000; // D (0x2000000000000010) 
    12'hae8 : errs =          63'b010000000000000000000000000000000000000000000000000000000100000; // D (0x2000000000000020) 
    12'hce9 : errs =          63'b010000000000000000000000000000000000000000000000000000001000000; // D (0x2000000000000040) 
    12'h0eb : errs =          63'b010000000000000000000000000000000000000000000000000000010000000; // D (0x2000000000000080) 
    12'hdd6 : errs =          63'b010000000000000000000000000000000000000000000000000000100000000; // D (0x2000000000000100) 
    12'h295 : errs =          63'b010000000000000000000000000000000000000000000000000001000000000; // D (0x2000000000000200) 
    12'h92a : errs =          63'b010000000000000000000000000000000000000000000000000010000000000; // D (0x2000000000000400) 
    12'hb6d : errs =          63'b010000000000000000000000000000000000000000000000000100000000000; // D (0x2000000000000800) 
    12'hfe3 : errs =          63'b010000000000000000000000000000000000000000000000001000000000000; // D (0x2000000000001000) 
    12'h6ff : errs =          63'b010000000000000000000000000000000000000000000000010000000000000; // D (0x2000000000002000) 
    12'h1fe : errs =          63'b010000000000000000000000000000000000000000000000100000000000000; // D (0x2000000000004000) 
    12'hffc : errs =          63'b010000000000000000000000000000000000000000000001000000000000000; // D (0x2000000000008000) 
    12'h6c1 : errs =          63'b010000000000000000000000000000000000000000000010000000000000000; // D (0x2000000000010000) 
    12'h182 : errs =          63'b010000000000000000000000000000000000000000000100000000000000000; // D (0x2000000000020000) 
    12'hf04 : errs =          63'b010000000000000000000000000000000000000000001000000000000000000; // D (0x2000000000040000) 
    12'h731 : errs =          63'b010000000000000000000000000000000000000000010000000000000000000; // D (0x2000000000080000) 
    12'h262 : errs =          63'b010000000000000000000000000000000000000000100000000000000000000; // D (0x2000000000100000) 
    12'h8c4 : errs =          63'b010000000000000000000000000000000000000001000000000000000000000; // D (0x2000000000200000) 
    12'h8b1 : errs =          63'b010000000000000000000000000000000000000010000000000000000000000; // D (0x2000000000400000) 
    12'h85b : errs =          63'b010000000000000000000000000000000000000100000000000000000000000; // D (0x2000000000800000) 
    12'h98f : errs =          63'b010000000000000000000000000000000000001000000000000000000000000; // D (0x2000000001000000) 
    12'ha27 : errs =          63'b010000000000000000000000000000000000010000000000000000000000000; // D (0x2000000002000000) 
    12'hd77 : errs =          63'b010000000000000000000000000000000000100000000000000000000000000; // D (0x2000000004000000) 
    12'h3d7 : errs =          63'b010000000000000000000000000000000001000000000000000000000000000; // D (0x2000000008000000) 
    12'hbae : errs =          63'b010000000000000000000000000000000010000000000000000000000000000; // D (0x2000000010000000) 
    12'he65 : errs =          63'b010000000000000000000000000000000100000000000000000000000000000; // D (0x2000000020000000) 
    12'h5f3 : errs =          63'b010000000000000000000000000000001000000000000000000000000000000; // D (0x2000000040000000) 
    12'h7e6 : errs =          63'b010000000000000000000000000000010000000000000000000000000000000; // D (0x2000000080000000) 
    12'h3cc : errs =          63'b010000000000000000000000000000100000000000000000000000000000000; // D (0x2000000100000000) 
    12'hb98 : errs =          63'b010000000000000000000000000001000000000000000000000000000000000; // D (0x2000000200000000) 
    12'he09 : errs =          63'b010000000000000000000000000010000000000000000000000000000000000; // D (0x2000000400000000) 
    12'h52b : errs =          63'b010000000000000000000000000100000000000000000000000000000000000; // D (0x2000000800000000) 
    12'h656 : errs =          63'b010000000000000000000000001000000000000000000000000000000000000; // D (0x2000001000000000) 
    12'h0ac : errs =          63'b010000000000000000000000010000000000000000000000000000000000000; // D (0x2000002000000000) 
    12'hd58 : errs =          63'b010000000000000000000000100000000000000000000000000000000000000; // D (0x2000004000000000) 
    12'h389 : errs =          63'b010000000000000000000001000000000000000000000000000000000000000; // D (0x2000008000000000) 
    12'hb12 : errs =          63'b010000000000000000000010000000000000000000000000000000000000000; // D (0x2000010000000000) 
    12'hf1d : errs =          63'b010000000000000000000100000000000000000000000000000000000000000; // D (0x2000020000000000) 
    12'h703 : errs =          63'b010000000000000000001000000000000000000000000000000000000000000; // D (0x2000040000000000) 
    12'h206 : errs =          63'b010000000000000000010000000000000000000000000000000000000000000; // D (0x2000080000000000) 
    12'h80c : errs =          63'b010000000000000000100000000000000000000000000000000000000000000; // D (0x2000100000000000) 
    12'h921 : errs =          63'b010000000000000001000000000000000000000000000000000000000000000; // D (0x2000200000000000) 
    12'hb7b : errs =          63'b010000000000000010000000000000000000000000000000000000000000000; // D (0x2000400000000000) 
    12'hfcf : errs =          63'b010000000000000100000000000000000000000000000000000000000000000; // D (0x2000800000000000) 
    12'h6a7 : errs =          63'b010000000000001000000000000000000000000000000000000000000000000; // D (0x2001000000000000) 
    12'h14e : errs =          63'b010000000000010000000000000000000000000000000000000000000000000; // D (0x2002000000000000) 
    12'he9c : errs =          63'b010000000000100000000000000000000000000000000000000000000000000; // D (0x2004000000000000) 
    12'h401 : errs =          63'b010000000001000000000000000000000000000000000000000000000000000; // D (0x2008000000000000) 
    12'h402 : errs =          63'b010000000010000000000000000000000000000000000000000000000000000; // D (0x2010000000000000) 
    12'h404 : errs =          63'b010000000100000000000000000000000000000000000000000000000000000; // D (0x2020000000000000) 
    12'h408 : errs =          63'b010000001000000000000000000000000000000000000000000000000000000; // D (0x2040000000000000) 
    12'h410 : errs =          63'b010000010000000000000000000000000000000000000000000000000000000; // D (0x2080000000000000) 
    12'h420 : errs =          63'b010000100000000000000000000000000000000000000000000000000000000; // D (0x2100000000000000) 
    12'h440 : errs =          63'b010001000000000000000000000000000000000000000000000000000000000; // D (0x2200000000000000) 
    12'h480 : errs =          63'b010010000000000000000000000000000000000000000000000000000000000; // D (0x2400000000000000) 
    12'h500 : errs =          63'b010100000000000000000000000000000000000000000000000000000000000; // D (0x2800000000000000) 
    12'h600 : errs =          63'b011000000000000000000000000000000000000000000000000000000000000; // D (0x3000000000000000) 
    12'h400 : errs =          63'b010000000000000000000000000000000000000000000000000000000000000; // S (0x2000000000000000) 
//    12'hc00 : errs =          63'b110000000000000000000000000000000000000000000000000000000000000; // D (0x6000000000000000) 
    12'hd39 : errs =          63'b100000000000000000000000000000000000000000000000000000000000001; // D (0x4000000000000001) 
    12'h272 : errs =          63'b100000000000000000000000000000000000000000000000000000000000010; // D (0x4000000000000002) 
    12'h9dd : errs =          63'b100000000000000000000000000000000000000000000000000000000000100; // D (0x4000000000000004) 
    12'hbba : errs =          63'b100000000000000000000000000000000000000000000000000000000001000; // D (0x4000000000000008) 
    12'hf74 : errs =          63'b100000000000000000000000000000000000000000000000000000000010000; // D (0x4000000000000010) 
    12'h6e8 : errs =          63'b100000000000000000000000000000000000000000000000000000000100000; // D (0x4000000000000020) 
    12'h0e9 : errs =          63'b100000000000000000000000000000000000000000000000000000001000000; // D (0x4000000000000040) 
    12'hceb : errs =          63'b100000000000000000000000000000000000000000000000000000010000000; // D (0x4000000000000080) 
    12'h1d6 : errs =          63'b100000000000000000000000000000000000000000000000000000100000000; // D (0x4000000000000100) 
    12'he95 : errs =          63'b100000000000000000000000000000000000000000000000000001000000000; // D (0x4000000000000200) 
    12'h52a : errs =          63'b100000000000000000000000000000000000000000000000000010000000000; // D (0x4000000000000400) 
    12'h76d : errs =          63'b100000000000000000000000000000000000000000000000000100000000000; // D (0x4000000000000800) 
    12'h3e3 : errs =          63'b100000000000000000000000000000000000000000000000001000000000000; // D (0x4000000000001000) 
    12'haff : errs =          63'b100000000000000000000000000000000000000000000000010000000000000; // D (0x4000000000002000) 
    12'hdfe : errs =          63'b100000000000000000000000000000000000000000000000100000000000000; // D (0x4000000000004000) 
    12'h3fc : errs =          63'b100000000000000000000000000000000000000000000001000000000000000; // D (0x4000000000008000) 
    12'hac1 : errs =          63'b100000000000000000000000000000000000000000000010000000000000000; // D (0x4000000000010000) 
    12'hd82 : errs =          63'b100000000000000000000000000000000000000000000100000000000000000; // D (0x4000000000020000) 
    12'h304 : errs =          63'b100000000000000000000000000000000000000000001000000000000000000; // D (0x4000000000040000) 
    12'hb31 : errs =          63'b100000000000000000000000000000000000000000010000000000000000000; // D (0x4000000000080000) 
    12'he62 : errs =          63'b100000000000000000000000000000000000000000100000000000000000000; // D (0x4000000000100000) 
    12'h4c4 : errs =          63'b100000000000000000000000000000000000000001000000000000000000000; // D (0x4000000000200000) 
    12'h4b1 : errs =          63'b100000000000000000000000000000000000000010000000000000000000000; // D (0x4000000000400000) 
    12'h45b : errs =          63'b100000000000000000000000000000000000000100000000000000000000000; // D (0x4000000000800000) 
    12'h58f : errs =          63'b100000000000000000000000000000000000001000000000000000000000000; // D (0x4000000001000000) 
    12'h627 : errs =          63'b100000000000000000000000000000000000010000000000000000000000000; // D (0x4000000002000000) 
    12'h177 : errs =          63'b100000000000000000000000000000000000100000000000000000000000000; // D (0x4000000004000000) 
    12'hfd7 : errs =          63'b100000000000000000000000000000000001000000000000000000000000000; // D (0x4000000008000000) 
    12'h7ae : errs =          63'b100000000000000000000000000000000010000000000000000000000000000; // D (0x4000000010000000) 
    12'h265 : errs =          63'b100000000000000000000000000000000100000000000000000000000000000; // D (0x4000000020000000) 
    12'h9f3 : errs =          63'b100000000000000000000000000000001000000000000000000000000000000; // D (0x4000000040000000) 
    12'hbe6 : errs =          63'b100000000000000000000000000000010000000000000000000000000000000; // D (0x4000000080000000) 
    12'hfcc : errs =          63'b100000000000000000000000000000100000000000000000000000000000000; // D (0x4000000100000000) 
    12'h798 : errs =          63'b100000000000000000000000000001000000000000000000000000000000000; // D (0x4000000200000000) 
    12'h209 : errs =          63'b100000000000000000000000000010000000000000000000000000000000000; // D (0x4000000400000000) 
    12'h92b : errs =          63'b100000000000000000000000000100000000000000000000000000000000000; // D (0x4000000800000000) 
    12'ha56 : errs =          63'b100000000000000000000000001000000000000000000000000000000000000; // D (0x4000001000000000) 
    12'hcac : errs =          63'b100000000000000000000000010000000000000000000000000000000000000; // D (0x4000002000000000) 
    12'h158 : errs =          63'b100000000000000000000000100000000000000000000000000000000000000; // D (0x4000004000000000) 
    12'hf89 : errs =          63'b100000000000000000000001000000000000000000000000000000000000000; // D (0x4000008000000000) 
    12'h712 : errs =          63'b100000000000000000000010000000000000000000000000000000000000000; // D (0x4000010000000000) 
    12'h31d : errs =          63'b100000000000000000000100000000000000000000000000000000000000000; // D (0x4000020000000000) 
    12'hb03 : errs =          63'b100000000000000000001000000000000000000000000000000000000000000; // D (0x4000040000000000) 
    12'he06 : errs =          63'b100000000000000000010000000000000000000000000000000000000000000; // D (0x4000080000000000) 
    12'h40c : errs =          63'b100000000000000000100000000000000000000000000000000000000000000; // D (0x4000100000000000) 
    12'h521 : errs =          63'b100000000000000001000000000000000000000000000000000000000000000; // D (0x4000200000000000) 
    12'h77b : errs =          63'b100000000000000010000000000000000000000000000000000000000000000; // D (0x4000400000000000) 
    12'h3cf : errs =          63'b100000000000000100000000000000000000000000000000000000000000000; // D (0x4000800000000000) 
    12'haa7 : errs =          63'b100000000000001000000000000000000000000000000000000000000000000; // D (0x4001000000000000) 
    12'hd4e : errs =          63'b100000000000010000000000000000000000000000000000000000000000000; // D (0x4002000000000000) 
    12'h29c : errs =          63'b100000000000100000000000000000000000000000000000000000000000000; // D (0x4004000000000000) 
    12'h801 : errs =          63'b100000000001000000000000000000000000000000000000000000000000000; // D (0x4008000000000000) 
    12'h802 : errs =          63'b100000000010000000000000000000000000000000000000000000000000000; // D (0x4010000000000000) 
    12'h804 : errs =          63'b100000000100000000000000000000000000000000000000000000000000000; // D (0x4020000000000000) 
    12'h808 : errs =          63'b100000001000000000000000000000000000000000000000000000000000000; // D (0x4040000000000000) 
    12'h810 : errs =          63'b100000010000000000000000000000000000000000000000000000000000000; // D (0x4080000000000000) 
    12'h820 : errs =          63'b100000100000000000000000000000000000000000000000000000000000000; // D (0x4100000000000000) 
    12'h840 : errs =          63'b100001000000000000000000000000000000000000000000000000000000000; // D (0x4200000000000000) 
    12'h880 : errs =          63'b100010000000000000000000000000000000000000000000000000000000000; // D (0x4400000000000000) 
    12'h900 : errs =          63'b100100000000000000000000000000000000000000000000000000000000000; // D (0x4800000000000000) 
    12'ha00 : errs =          63'b101000000000000000000000000000000000000000000000000000000000000; // D (0x5000000000000000) 
    12'hc00 : errs =          63'b110000000000000000000000000000000000000000000000000000000000000; // D (0x6000000000000000) 
    12'h800 : errs =          63'b100000000000000000000000000000000000000000000000000000000000000; // S (0x4000000000000000) 

default : errs = {(31){1'b0}};     
 endcase	

// Num of errs. =        3969. Single =          63. Double =        3906

 fn_err_pat_dcd_gf6_rom = errs; 
 
end						
endfunction // fn_err_pat_dcd_gf6_rom			
